/*
* Copyright 2018-2022 F4PGA Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0
*/

/*
 * Generated by harness_gen.py
 * From: simpleuart.v
 */
module top(input wire clk, input wire stb, input wire di, output wire do);
    localparam integer DIN_N = 72;
    localparam integer DOUT_N = 66;

    reg [DIN_N-1:0] din;
    wire [DOUT_N-1:0] dout;

    reg [DIN_N-1:0] din_shr;
    reg [DOUT_N-1:0] dout_shr;

    always @(posedge clk) begin
        din_shr <= {din_shr, di};
        dout_shr <= {dout_shr, din_shr[DIN_N-1]};
        if (stb) begin
            din <= din_shr;
            dout_shr <= dout;
        end
    end

    assign do = dout_shr[DOUT_N-1];
    simpleuart dut(
            .clk(clk),
            .resetn(din[0]),
            .ser_tx(dout[0]),
            .ser_rx(din[1]),
            .reg_div_we(din[5:2]),
            .reg_div_di(din[37:6]),
            .reg_div_do(dout[32:1]),
            .reg_dat_we(din[38]),
            .reg_dat_re(din[39]),
            .reg_dat_di(din[71:40]),
            .reg_dat_do(dout[64:33]),
            .reg_dat_wait(dout[65])
            );
endmodule
