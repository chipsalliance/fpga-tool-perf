/* Machine-generated using LiteX gen */
module top(
	output reg serial_tx,
	input serial_rx,
	input clk50,
	output [13:0] ddram_a,
	output [2:0] ddram_ba,
	output ddram_ras_n,
	output ddram_cas_n,
	output ddram_we_n,
	output [3:0] ddram_dm,
	inout [31:0] ddram_dq,
	output [3:0] ddram_dqs_p,
	output [3:0] ddram_dqs_n,
	output ddram_clk_p,
	output ddram_clk_n,
	output ddram_cke,
	output ddram_odt,
	output ddram_reset_n,
	output ddram_cs_n,
	output fpga_led00,
	output fpga_led10,
	input hdmi_in0_clk_p,
	input hdmi_in0_clk_n,
	input hdmi_in0_data0_p,
	input hdmi_in0_data0_n,
	input hdmi_in0_data1_p,
	input hdmi_in0_data1_n,
	input hdmi_in0_data2_p,
	input hdmi_in0_data2_n,
	input hdmi_in0_scl,
	inout hdmi_in0_sda,
	input hdmi_in0_hpd_notif,
	output hdmi_out0_clk_p,
	output hdmi_out0_clk_n,
	output hdmi_out0_data0_p,
	output hdmi_out0_data0_n,
	output hdmi_out0_data1_p,
	output hdmi_out0_data1_n,
	output hdmi_out0_data2_p,
	output hdmi_out0_data2_n,
	output hdmi_sda_over_up,
	output hdmi_sda_over_dn,
	input hdmi_in1_clk_p,
	input hdmi_in1_clk_n,
	input hdmi_in1_data0_p,
	input hdmi_in1_data0_n,
	input hdmi_in1_data1_p,
	input hdmi_in1_data1_n,
	input hdmi_in1_data2_p,
	input hdmi_in1_data2_n,
	input hdmi_in1_scl,
	inout hdmi_in1_sda,
	output hpd_en,
	output fpga_led20,
	output fpga_led30,
	output fpga_led50,
	output rmii_eth_clocks_ref_clk,
	output rmii_eth_rst_n,
	input [1:0] rmii_eth_rx_data,
	input rmii_eth_crs_dv,
	output reg rmii_eth_tx_en,
	output reg [1:0] rmii_eth_tx_data,
	output rmii_eth_mdc,
	inout rmii_eth_mdio,
	input rmii_eth_rx_er,
	input rmii_eth_int_n,
	output reg fpga_led40
);

wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_reset_reset_re;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_reset_reset_r;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_reset_reset_w = 1'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full = 32'd305419896;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_re = 1'd0;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors_status;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_reset;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_error;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors = 32'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_reset;
wire [29:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_adr;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_dat_w;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_dat_r;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_sel;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_cyc;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_stb;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_ack;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_we;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_cti;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_bte;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_err = 1'd0;
wire [29:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_adr;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_dat_w;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_dat_r;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_sel;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_cyc;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_stb;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_ack;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_we;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_cti;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_bte;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_err = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_err = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_d_err = 1'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_interrupt = 32'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_reset = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_cpu_reset = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_wr = 1'd0;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_address = 8'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_data = 32'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_o_cmd_ready;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_o_rsp_data;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_o_resetOut;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_reset_debug_logic = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_complete = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_in_progress = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_wait_for_ack = 1'd0;
wire [29:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_adr;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_dat_w;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_dat_r = 32'd0;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_sel;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_cyc;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_stb;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_ack = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_we;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_cti;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_bte;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_err = 1'd0;
wire [29:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_adr;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_dat_w;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_dat_r;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_sel;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_cyc;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_stb;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_ack = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_we;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_cti;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_bte;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_err = 1'd0;
wire [12:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_adr;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_dat_r;
wire [29:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_adr;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_dat_w;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_dat_r;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_sel;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_cyc;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_stb;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_ack = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_we;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_cti;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_bte;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_err = 1'd0;
wire [11:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_adr;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_dat_r;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_we = 4'd0;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_dat_w;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr = 14'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we = 1'd0;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w = 8'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_r;
wire [29:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_adr;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_dat_w;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_dat_r = 32'd0;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_sel;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_cyc;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_stb;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_ack = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_we;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_cti;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_bte;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_err = 1'd0;
reg [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_counter = 2'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full = 32'd4947802;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_re = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_valid;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_ready = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_first;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_last;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_payload_data;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_uart_clk_txen = 1'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_phase_accumulator_tx = 32'd0;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_reg = 8'd0;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_bitcount = 4'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_busy = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_ready;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_first = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_payload_data = 8'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_uart_clk_rxen = 1'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_phase_accumulator_rx = 32'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_r = 1'd0;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_reg = 8'd0;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_bitcount = 4'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_busy = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxtx_re;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxtx_r;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxtx_w;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_txfull_status;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxempty_status;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_irq;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_status;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_pending = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_trigger;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_clear = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_old_trigger = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_status;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_pending = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_trigger;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_clear = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_old_trigger = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_status_re;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_status_r;
reg [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_status_w = 2'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_re;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_r;
reg [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_w = 2'd0;
reg [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_storage_full = 2'd0;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_storage;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_re = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_ready;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_first = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_last = 1'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_payload_data;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_first;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_last;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_payload_data;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_re;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_readable = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_we;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_writable;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_re;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_readable;
wire [9:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_din;
wire [9:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_dout;
reg [4:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level0 = 5'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_replace = 1'd0;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_produce = 4'd0;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_consume = 4'd0;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_adr = 4'd0;
wire [9:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_we;
wire [9:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_dat_w;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_do_read;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_rdport_adr;
wire [9:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_rdport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_rdport_re;
wire [4:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level1;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_in_payload_data;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_in_first;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_in_last;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_out_payload_data;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_out_first;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_out_last;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_ready;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_first;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_last;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_payload_data;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_first;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_last;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_payload_data;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_re;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_readable = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_we;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_writable;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_re;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_readable;
wire [9:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_din;
wire [9:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_dout;
reg [4:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level0 = 5'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_replace = 1'd0;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_produce = 4'd0;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_consume = 4'd0;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_adr = 4'd0;
wire [9:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_we;
wire [9:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_dat_w;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_do_read;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_rdport_adr;
wire [9:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_rdport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_rdport_re;
wire [4:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level1;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_in_payload_data;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_in_first;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_in_last;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_out_payload_data;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_out_first;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_out_last;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_reset;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full = 32'd0;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_re = 1'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full = 32'd0;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_re = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_storage_full = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_storage;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_re = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_update_value_re;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_update_value_r;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_update_value_w = 1'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value_status = 32'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_irq;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_status;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_pending = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_trigger;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_clear = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_old_trigger = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_status_re;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_status_r;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_status_w;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_pending_re;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_pending_r;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_pending_w;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_storage_full = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_storage;
reg soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_re = 1'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value = 32'd0;
wire [29:0] soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_w;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r = 32'd0;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_sel;
wire soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_cyc;
wire soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_stb;
reg soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_ack = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_we;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_cti;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_bte;
reg soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_err = 1'd0;
(* dont_touch = "true" *) wire sys_clk;
wire sys_rst;
wire sys4x_clk;
wire sys4x_dqs_clk;
wire clk200_clk;
wire clk200_rst;
wire eth_clk;
wire eth_rst;
reg soc_videooverlaysoc_videooverlaysoc_crg_rst = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_crg_pll_locked;
wire soc_videooverlaysoc_videooverlaysoc_crg_pll_fb;
wire soc_videooverlaysoc_videooverlaysoc_crg_pll_sys;
wire soc_videooverlaysoc_videooverlaysoc_crg_pll_sys4x;
wire soc_videooverlaysoc_videooverlaysoc_crg_pll_sys4x_dqs;
wire soc_videooverlaysoc_videooverlaysoc_crg_pll_clk200;
wire soc_videooverlaysoc_videooverlaysoc_crg_pll_clk50;
wire soc_videooverlaysoc_videooverlaysoc_crg_pll_fb_bufg;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_crg_reset_counter = 4'd15;
reg soc_videooverlaysoc_videooverlaysoc_crg_ic_reset = 1'd1;
reg [11:0] soc_videooverlaysoc_videooverlaysoc_temperature_status = 12'd0;
reg [11:0] soc_videooverlaysoc_videooverlaysoc_vccint_status = 12'd0;
reg [11:0] soc_videooverlaysoc_videooverlaysoc_vccaux_status = 12'd0;
reg [11:0] soc_videooverlaysoc_videooverlaysoc_vccbram_status = 12'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_alarm;
wire soc_videooverlaysoc_videooverlaysoc_ot;
wire soc_videooverlaysoc_videooverlaysoc_busy;
wire [6:0] soc_videooverlaysoc_videooverlaysoc_channel;
wire soc_videooverlaysoc_videooverlaysoc_eoc;
wire soc_videooverlaysoc_videooverlaysoc_eos;
wire [15:0] soc_videooverlaysoc_videooverlaysoc_data;
wire soc_videooverlaysoc_videooverlaysoc_drdy;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_half_sys8x_taps_storage_full = 4'd8;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_half_sys8x_taps_storage;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_half_sys8x_taps_re = 1'd0;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage_full = 4'd0;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_re = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_r;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_w = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_r;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_w = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_r;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_w = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_r;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_w = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_bank;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cas_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cs_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_ras_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_we_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cke;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_odt;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_reset_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_act_n;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata_valid = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_bank;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cas_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cs_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_ras_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_we_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cke;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_odt;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_reset_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_act_n;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata_valid = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_bank;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cas_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cs_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_ras_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_we_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cke;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_odt;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_reset_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_act_n;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata_valid = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_bank;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cas_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cs_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_ras_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_we_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cke;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_odt;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_reset_n;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_act_n;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_sd_clk_se;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dqs = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_preamble;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_postamble;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern = 8'd85;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay1;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t1;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy1;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay2;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t2;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy2;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay3;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t3;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy3;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay1;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay1;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed1;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t1;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data1;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay2;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay2;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed2;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t2;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data2;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay3;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay3;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed3;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t3;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data3;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay4;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay4;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed4;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t4;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data4;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay5;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay5;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed5;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t5;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data5;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay6;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay6;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed6;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t6;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data6;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay7;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay7;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed7;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t7;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data7;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay8;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay8;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed8;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t8;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data8;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay9;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay9;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed9;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t9;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data9;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay10;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay10;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed10;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t10;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data10;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay11;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay11;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed11;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t11;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data11;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay12;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay12;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed12;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t12;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data12;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay13;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay13;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed13;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t13;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data13;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay14;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay14;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed14;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t14;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data14;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay15;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay15;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed15;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t15;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data15;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay16;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay16;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed16;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t16;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data16;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay17;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay17;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed17;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t17;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data17;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay18;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay18;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed18;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t18;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data18;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay19;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay19;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed19;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t19;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data19;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay20;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay20;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed20;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t20;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data20;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay21;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay21;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed21;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t21;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data21;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay22;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay22;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed22;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t22;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data22;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay23;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay23;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed23;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t23;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data23;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay24;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay24;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed24;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t24;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data24;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay25;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay25;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed25;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t25;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data25;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay26;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay26;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed26;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t26;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data26;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay27;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay27;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed27;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t27;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data27;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay28;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay28;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed28;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t28;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data28;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay29;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay29;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed29;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t29;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data29;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay30;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay30;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed30;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t30;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data30;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r = 16'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay31;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay31;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed31;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t31;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data31;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_i;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o = 8'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_value = 3'd0;
reg [15:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r = 16'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en0 = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en1 = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en2 = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en3 = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en4 = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en5 = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en6 = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en7 = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en = 4'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_bank;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_we_n = 1'd1;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_reset_n;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_act_n = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata_valid = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_bank;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_we_n = 1'd1;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_reset_n;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_act_n = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata_valid = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_bank;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_we_n = 1'd1;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_reset_n;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_act_n = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata_valid = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_bank;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_we_n = 1'd1;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_reset_n;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_act_n = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata_valid = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_bank;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_cas_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_cs_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_ras_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_we_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_reset_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_act_n;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata_valid = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_bank;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_cas_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_cs_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_ras_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_we_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_reset_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_act_n;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata_valid = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_bank;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_cas_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_cs_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_ras_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_we_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_reset_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_act_n;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata_valid = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_address;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_bank;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_cas_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_cs_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_ras_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_we_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_reset_n;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_act_n;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_wrdata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_wrdata_en;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_wrdata_mask;
wire soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata_en;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata_valid = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_address = 14'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_bank = 3'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_we_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cke = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_odt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_reset_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_act_n = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata_en = 1'd0;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata_mask = 8'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata_en = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata_valid;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_address = 14'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_bank = 3'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_we_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cke = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_odt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_reset_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_act_n = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata_en = 1'd0;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata_mask = 8'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata_en = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata_valid;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_address = 14'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_bank = 3'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_we_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cke = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_odt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_reset_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_act_n = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata_en = 1'd0;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata_mask = 8'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata_en = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata_valid;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_address = 14'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_bank = 3'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_we_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cke = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_odt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_reset_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_act_n = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata = 64'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata_en = 1'd0;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata_mask = 8'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata_en = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata_valid;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_storage_full = 4'd0;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_re = 1'd0;
reg [5:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage_full = 6'd0;
wire [5:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_re = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_issue_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_issue_r;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_issue_w = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_storage_full = 14'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_re = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_storage_full = 3'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_re = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full = 64'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_re = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status = 64'd0;
reg [5:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage_full = 6'd0;
wire [5:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_re = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_issue_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_issue_r;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_issue_w = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_storage_full = 14'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_re = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_storage_full = 3'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_re = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full = 64'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_re = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status = 64'd0;
reg [5:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage_full = 6'd0;
wire [5:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_re = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_issue_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_issue_r;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_issue_w = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_storage_full = 14'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_re = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_storage_full = 3'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_re = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full = 64'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_re = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status = 64'd0;
reg [5:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage_full = 6'd0;
wire [5:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_re = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_issue_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_issue_r;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_issue_w = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_storage_full = 14'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_re = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_storage_full = 3'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_re = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full = 64'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage;
reg soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_re = 1'd0;
reg [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status = 64'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_address = 14'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_bank = 3'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_we_n = 1'd1;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_reset_n;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_act_n = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_wrdata;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_wrdata_en = 1'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_wrdata_mask;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_rddata_en = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_rddata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_rddata_valid;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_address = 14'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_bank = 3'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_we_n = 1'd1;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_reset_n;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_act_n = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_wrdata;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_wrdata_en = 1'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_wrdata_mask;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_rddata_en = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_rddata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_rddata_valid;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_address = 14'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_bank = 3'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_we_n = 1'd1;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_reset_n;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_act_n = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_wrdata;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_wrdata_en = 1'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_wrdata_mask;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_rddata_en = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_rddata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_rddata_valid;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_address = 14'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_bank = 3'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cas_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cs_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_ras_n = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_we_n = 1'd1;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cke;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_odt;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_reset_n;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_act_n = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_wrdata;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_wrdata_en = 1'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_wrdata_mask;
reg soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_rddata_en = 1'd0;
wire [63:0] soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_rddata;
wire soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_rddata_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_wdata_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_rdata_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_wdata_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_rdata_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_wdata_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_rdata_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_wdata_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_rdata_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_wdata_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_rdata_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_wdata_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_rdata_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_wdata_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_rdata_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_wdata_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_rdata_valid;
reg [255:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata = 256'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata_we = 32'd0;
wire [255:0] soc_videooverlaysoc_videooverlaysoc_sdram_interface_rdata;
reg soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_cmd_last = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_a = 14'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ba = 3'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_we = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_is_read = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_is_write = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_seq_start = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_seq_done = 1'd0;
reg [4:0] soc_videooverlaysoc_videooverlaysoc_sdram_counter = 5'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_wait;
wire soc_videooverlaysoc_videooverlaysoc_sdram_done;
reg [9:0] soc_videooverlaysoc_videooverlaysoc_sdram_count = 10'd782;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_lock;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_wdata_ready = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_rdata_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_refresh_req;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_refresh_gnt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_a = 14'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ba;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_we = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_cmd = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_read = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_write = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_auto_precharge = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_ready;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_first = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_last = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_we;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_readable;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_din;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_dout;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_level = 4'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_we;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_dat_w;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_do_read;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_rdport_adr;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_rdport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_last;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_addr = 21'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_pipe_ce;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_busy;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_valid_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_first_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_last_n = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row = 14'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_opened = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_hit;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_open = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_close = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_col_n_addr_sel = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_lock;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_wdata_ready = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_rdata_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_refresh_req;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_refresh_gnt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_a = 14'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ba;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_we = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_cmd = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_read = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_write = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_auto_precharge = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_ready;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_first = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_last = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_we;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_readable;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_din;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_dout;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_level = 4'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_we;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_dat_w;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_do_read;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_rdport_adr;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_rdport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_last;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_addr = 21'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_pipe_ce;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_busy;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_valid_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_first_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_last_n = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row = 14'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_opened = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_hit;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_open = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_close = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_col_n_addr_sel = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_lock;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_wdata_ready = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_rdata_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_refresh_req;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_refresh_gnt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_a = 14'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ba;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_we = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_cmd = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_read = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_write = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_auto_precharge = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_ready;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_first = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_last = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_we;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_readable;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_din;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_dout;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_level = 4'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_we;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_dat_w;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_do_read;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_rdport_adr;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_rdport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_last;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_addr = 21'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_pipe_ce;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_busy;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_valid_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_first_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_last_n = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row = 14'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_opened = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_hit;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_open = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_close = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_col_n_addr_sel = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_lock;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_wdata_ready = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_rdata_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_refresh_req;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_refresh_gnt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_a = 14'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ba;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_we = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_cmd = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_read = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_write = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_auto_precharge = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_ready;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_first = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_last = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_we;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_readable;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_din;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_dout;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_level = 4'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_we;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_dat_w;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_do_read;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_rdport_adr;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_rdport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_last;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_addr = 21'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_pipe_ce;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_busy;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_valid_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_first_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_last_n = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row = 14'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_opened = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_hit;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_open = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_close = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_col_n_addr_sel = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_lock;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_wdata_ready = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_rdata_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_refresh_req;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_refresh_gnt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_a = 14'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ba;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_we = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_cmd = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_read = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_write = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_auto_precharge = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_ready;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_first = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_last = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_we;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_readable;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_din;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_dout;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_level = 4'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_we;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_dat_w;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_do_read;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_rdport_adr;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_rdport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_last;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_addr = 21'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_pipe_ce;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_busy;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_valid_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_first_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_last_n = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row = 14'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_opened = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_hit;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_open = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_close = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_col_n_addr_sel = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_lock;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_wdata_ready = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_rdata_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_refresh_req;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_refresh_gnt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_a = 14'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ba;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_we = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_cmd = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_read = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_write = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_auto_precharge = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_ready;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_first = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_last = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_we;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_readable;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_din;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_dout;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_level = 4'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_we;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_dat_w;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_do_read;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_rdport_adr;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_rdport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_last;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_addr = 21'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_pipe_ce;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_busy;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_valid_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_first_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_last_n = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row = 14'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_opened = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_hit;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_open = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_close = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_col_n_addr_sel = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_lock;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_wdata_ready = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_rdata_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_refresh_req;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_refresh_gnt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_a = 14'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ba;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_we = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_cmd = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_read = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_write = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_auto_precharge = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_ready;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_first = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_last = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_we;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_readable;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_din;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_dout;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_level = 4'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_we;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_dat_w;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_do_read;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_rdport_adr;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_rdport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_last;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_addr = 21'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_pipe_ce;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_busy;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_valid_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_first_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_last_n = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row = 14'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_opened = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_hit;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_open = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_close = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_col_n_addr_sel = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_lock;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_wdata_ready = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_rdata_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_refresh_req;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_refresh_gnt = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_a = 14'd0;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ba;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_we = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_cmd = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_read = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_write = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_auto_precharge = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_ready;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_first = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_last = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_we;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_readable;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_din;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_dout;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_level = 4'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_we;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_dat_w;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_do_read;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_rdport_adr;
wire [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_rdport_dat_r;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_last;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_payload_we;
wire [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_payload_addr;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_valid;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_ready;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_first;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_last;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_addr = 21'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_pipe_ce;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_busy;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_valid_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_first_n = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_last_n = 1'd0;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row = 14'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_opened = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_hit;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_open = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_close = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_col_n_addr_sel = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_ras_allowed;
wire soc_videooverlaysoc_videooverlaysoc_sdram_cas_allowed;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_reads = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_writes = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_cmds = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_a;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ba;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_cmd;
wire soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_read;
wire soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_write;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids = 8'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_ce;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_cmds = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_activates = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready = 1'd0;
wire [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_a;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ba;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_cas = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ras = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_we = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_cmd;
wire soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_read;
wire soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_write;
reg [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids = 8'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_ce;
reg [13:0] soc_videooverlaysoc_videooverlaysoc_sdram_nop_a = 14'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_nop_ba = 3'd0;
reg [1:0] soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0 = 2'd0;
reg [1:0] soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1 = 2'd0;
reg [1:0] soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2 = 2'd0;
reg [1:0] soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3 = 2'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_steerer0 = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_steerer1 = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_steerer2 = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_steerer3 = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_steerer4 = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_steerer5 = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_steerer6 = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_steerer7 = 1'd1;
wire soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_ready = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_count = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_ready = 1'd1;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_count;
reg [4:0] soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_window = 5'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_ready = 1'd1;
reg soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_count = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_valid;
(* dont_touch = "true" *) reg soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_ready = 1'd1;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_count = 3'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_read_available;
wire soc_videooverlaysoc_videooverlaysoc_sdram_write_available;
reg soc_videooverlaysoc_videooverlaysoc_sdram_en0 = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_max_time0;
reg [4:0] soc_videooverlaysoc_videooverlaysoc_sdram_time0 = 5'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_en1 = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_max_time1;
reg [3:0] soc_videooverlaysoc_videooverlaysoc_sdram_time1 = 4'd0;
wire soc_videooverlaysoc_videooverlaysoc_sdram_go_to_refresh;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_update_re;
wire soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_update_r;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_update_w = 1'd0;
reg [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads_status = 24'd0;
reg [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites_status = 24'd0;
reg [8:0] soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_data_width_status = 9'd256;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_valid = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_ready = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_is_read = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_is_write = 1'd0;
reg [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_counter = 24'd0;
reg soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_period = 1'd0;
reg [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads = 24'd0;
reg [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites = 24'd0;
reg [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads_r = 24'd0;
reg [23:0] soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites_r = 24'd0;
wire [29:0] soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_adr;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_dat_w;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_dat_r;
wire [3:0] soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_sel;
wire soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_cyc;
wire soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_stb;
wire soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_ack;
wire soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_we;
wire [2:0] soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_cti;
wire [1:0] soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_bte;
wire soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_err;
reg soc_videooverlaysoc_videooverlaysoc_port_cmd_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_port_cmd_ready;
reg soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we = 1'd0;
reg [23:0] soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr = 24'd0;
reg soc_videooverlaysoc_videooverlaysoc_port_wdata_valid = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_port_wdata_ready;
reg [255:0] soc_videooverlaysoc_videooverlaysoc_port_wdata_payload_data = 256'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_port_wdata_payload_we = 32'd0;
wire soc_videooverlaysoc_videooverlaysoc_port_rdata_valid;
reg soc_videooverlaysoc_videooverlaysoc_port_rdata_ready = 1'd0;
wire [255:0] soc_videooverlaysoc_videooverlaysoc_port_rdata_payload_data;
wire [29:0] soc_videooverlaysoc_videooverlaysoc_adr;
wire [255:0] soc_videooverlaysoc_videooverlaysoc_dat_w;
reg [255:0] soc_videooverlaysoc_videooverlaysoc_dat_r = 256'd0;
wire [31:0] soc_videooverlaysoc_videooverlaysoc_sel;
reg soc_videooverlaysoc_videooverlaysoc_cyc = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_stb = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_ack = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_we = 1'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_data_port_adr;
wire [255:0] soc_videooverlaysoc_videooverlaysoc_data_port_dat_r;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_data_port_we = 32'd0;
reg [255:0] soc_videooverlaysoc_videooverlaysoc_data_port_dat_w = 256'd0;
reg soc_videooverlaysoc_videooverlaysoc_write_from_slave = 1'd0;
reg [2:0] soc_videooverlaysoc_videooverlaysoc_adr_offset_r = 3'd0;
wire [7:0] soc_videooverlaysoc_videooverlaysoc_tag_port_adr;
wire [25:0] soc_videooverlaysoc_videooverlaysoc_tag_port_dat_r;
reg soc_videooverlaysoc_videooverlaysoc_tag_port_we = 1'd0;
wire [25:0] soc_videooverlaysoc_videooverlaysoc_tag_port_dat_w;
wire [24:0] soc_videooverlaysoc_videooverlaysoc_tag_do_tag;
wire soc_videooverlaysoc_videooverlaysoc_tag_do_dirty;
wire [24:0] soc_videooverlaysoc_videooverlaysoc_tag_di_tag;
reg soc_videooverlaysoc_videooverlaysoc_tag_di_dirty = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_word_clr = 1'd0;
reg soc_videooverlaysoc_videooverlaysoc_word_inc = 1'd0;
wire soc_videooverlaysoc_videooverlaysoc_sys_led;
reg soc_videooverlaysoc_videooverlaysoc_pcie_led = 1'd0;
reg [31:0] soc_videooverlaysoc_videooverlaysoc_sys_counter = 32'd0;
wire soc_videooverlaysoc_hdmi_in0_freq_clk0;
wire [31:0] soc_videooverlaysoc_hdmi_in0_freq_status;
wire hdmi_in0_freq_fmeter_clk;
wire soc_videooverlaysoc_hdmi_in0_freq_period_done;
reg [31:0] soc_videooverlaysoc_hdmi_in0_freq_period_counter = 32'd0;
wire soc_videooverlaysoc_hdmi_in0_freq_ce;
reg [5:0] soc_videooverlaysoc_hdmi_in0_freq_q = 6'd0;
wire [5:0] soc_videooverlaysoc_hdmi_in0_freq_q_next;
reg [5:0] soc_videooverlaysoc_hdmi_in0_freq_q_binary = 6'd0;
reg [5:0] soc_videooverlaysoc_hdmi_in0_freq_q_next_binary = 6'd0;
wire [5:0] soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_i;
reg [5:0] soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o = 6'd0;
reg [5:0] soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb = 6'd0;
wire soc_videooverlaysoc_hdmi_in0_freq_sampler_latch;
wire [5:0] soc_videooverlaysoc_hdmi_in0_freq_sampler_i;
reg [31:0] soc_videooverlaysoc_hdmi_in0_freq_sampler_o = 32'd0;
wire [5:0] soc_videooverlaysoc_hdmi_in0_freq_sampler_inc;
reg [31:0] soc_videooverlaysoc_hdmi_in0_freq_sampler_counter = 32'd0;
reg [5:0] soc_videooverlaysoc_hdmi_in0_freq_sampler_i_d = 6'd0;
wire soc_videooverlaysoc_hdmi_in0_edid_status;
reg soc_videooverlaysoc_hdmi_in0_edid_storage_full = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_edid_storage;
reg soc_videooverlaysoc_hdmi_in0_edid_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_edid_hpd_notif_n;
wire soc_videooverlaysoc_hdmi_in0_edid_scl_raw;
reg soc_videooverlaysoc_hdmi_in0_edid_sda_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_edid_sda_raw;
reg soc_videooverlaysoc_hdmi_in0_edid_sda_drv = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_sda_drv_reg = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_edid_sda_i_async;
wire soc_videooverlaysoc_hdmi_in0_edid_sda_o;
reg soc_videooverlaysoc_hdmi_in0_edid_scl_i = 1'd0;
reg [5:0] soc_videooverlaysoc_hdmi_in0_edid_samp_count = 6'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_samp_carry = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_scl_r = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_sda_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_edid_scl_rising;
wire soc_videooverlaysoc_hdmi_in0_edid_sda_rising;
wire soc_videooverlaysoc_hdmi_in0_edid_sda_falling;
wire soc_videooverlaysoc_hdmi_in0_edid_start;
reg [7:0] soc_videooverlaysoc_hdmi_in0_edid_din = 8'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_edid_counter = 4'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_is_read = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_update_is_read = 1'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_edid_offset_counter = 8'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_oc_load = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_oc_inc = 1'd0;
wire [7:0] soc_videooverlaysoc_hdmi_in0_edid_adr;
wire [7:0] soc_videooverlaysoc_hdmi_in0_edid_dat_r;
reg soc_videooverlaysoc_hdmi_in0_edid_data_bit = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_zero_drv = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_data_drv = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_data_drv_en = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_edid_data_drv_stop = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_mmcm_reset_storage_full = 1'd1;
wire soc_videooverlaysoc_hdmi_in0_mmcm_reset_storage;
reg soc_videooverlaysoc_hdmi_in0_mmcm_reset_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_locked_status;
wire soc_videooverlaysoc_hdmi_in0_mmcm_read_re;
wire soc_videooverlaysoc_hdmi_in0_mmcm_read_r;
reg soc_videooverlaysoc_hdmi_in0_mmcm_read_w = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_mmcm_write_re;
wire soc_videooverlaysoc_hdmi_in0_mmcm_write_r;
reg soc_videooverlaysoc_hdmi_in0_mmcm_write_w = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_mmcm_drdy_status = 1'd0;
reg [6:0] soc_videooverlaysoc_hdmi_in0_mmcm_adr_storage_full = 7'd0;
wire [6:0] soc_videooverlaysoc_hdmi_in0_mmcm_adr_storage;
reg soc_videooverlaysoc_hdmi_in0_mmcm_adr_re = 1'd0;
reg [15:0] soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage_full = 16'd0;
wire [15:0] soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage;
reg soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_re = 1'd0;
wire [15:0] soc_videooverlaysoc_hdmi_in0_mmcm_dat_r_status;
wire soc_videooverlaysoc_hdmi_in0_locked;
wire hdmi_in0_pix_clk;
wire hdmi_in0_pix_rst;
wire hdmi_in0_pix1p25x_clk;
wire hdmi_in0_pix1p25x_rst;
wire hdmi_in0_pix5x_clk;
wire soc_videooverlaysoc_hdmi_in0_mmcm_write_o_re;
wire soc_videooverlaysoc_hdmi_in0_mmcm_write_o_r;
reg soc_videooverlaysoc_hdmi_in0_mmcm_write_o_w = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_mmcm_read_o_re;
wire soc_videooverlaysoc_hdmi_in0_mmcm_read_o_r;
reg soc_videooverlaysoc_hdmi_in0_mmcm_read_o_w = 1'd0;
wire [15:0] soc_videooverlaysoc_hdmi_in0_mmcm_dat_o_r_status;
reg soc_videooverlaysoc_hdmi_in0_mmcm_drdy_o_status = 1'd0;
wire pix_o_clk;
wire pix_o_rst;
wire pix5x_o_clk;
wire soc_videooverlaysoc_hdmi_in0_clk_input;
wire soc_videooverlaysoc_hdmi_in0_clk_input_bufr;
wire soc_videooverlaysoc_hdmi_in0_mmcm_fb;
wire soc_videooverlaysoc_hdmi_in0_mmcm_locked;
wire soc_videooverlaysoc_hdmi_in0_mmcm_clk0;
wire soc_videooverlaysoc_hdmi_in0_mmcm_clk1;
wire soc_videooverlaysoc_hdmi_in0_mmcm_clk2;
wire soc_videooverlaysoc_hdmi_in0_mmcm_drdy;
wire soc_videooverlaysoc_hdmi_in0_mmcm_fb_o;
wire soc_videooverlaysoc_hdmi_in0_mmcm_fb2_o;
wire soc_videooverlaysoc_hdmi_in0_mmcm_locked_o;
wire soc_videooverlaysoc_hdmi_in0_mmcm_clk0_o;
wire soc_videooverlaysoc_hdmi_in0_mmcm_clk2_o;
wire soc_videooverlaysoc_hdmi_in0_mmcm_drdy_o;
wire [9:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_d;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_re;
wire [4:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_r;
reg [4:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_w = 5'd0;
wire [1:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_status;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_phase_reset_re;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_phase_reset_r;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_phase_reset_w = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_i_nodelay;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_i_nodelay;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_rst;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_master_inc;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_master_ce;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_slave_inc;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_slave_ce;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_q;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_d;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_q;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_d;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
reg [9:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_o = 10'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst_write = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst_read = 1'd0;
wire hdmi_in0_data0_cap_write_clk;
wire hdmi_in0_data0_cap_write_rst;
wire hdmi_in0_data0_cap_read_clk;
wire hdmi_in0_data0_cap_read_rst;
reg [79:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr = 80'd0;
reg [79:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_rd = 80'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_wrpointer = 4'd5;
reg [2:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rdpointer = 3'd0;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_mdata;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_sdata;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_inc;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_dec;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_transition;
reg [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_mdata_d = 8'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture0_lateness = 8'd128;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_too_late;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_too_early;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_reset_lateness;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_charsync0_raw_data;
reg soc_videooverlaysoc_hdmi_in0_charsync0_synced = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in0_charsync0_data = 10'd0;
wire soc_videooverlaysoc_hdmi_in0_charsync0_char_synced_status;
wire [3:0] soc_videooverlaysoc_hdmi_in0_charsync0_ctl_pos_status;
reg [9:0] soc_videooverlaysoc_hdmi_in0_charsync0_raw_data1 = 10'd0;
wire [19:0] soc_videooverlaysoc_hdmi_in0_charsync0_raw;
reg soc_videooverlaysoc_hdmi_in0_charsync0_found_control = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_charsync0_control_position = 4'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in0_charsync0_control_counter = 3'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_charsync0_previous_control_position = 4'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_charsync0_word_sel = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_wer0_data;
wire soc_videooverlaysoc_hdmi_in0_wer0_update_re;
wire soc_videooverlaysoc_hdmi_in0_wer0_update_r;
reg soc_videooverlaysoc_hdmi_in0_wer0_update_w = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer0_status = 24'd0;
reg [8:0] soc_videooverlaysoc_hdmi_in0_wer0_data_r = 9'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_wer0_transitions = 8'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_wer0_transition_count = 4'd0;
reg soc_videooverlaysoc_hdmi_in0_wer0_is_control = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_wer0_is_error = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer0_period_counter = 24'd0;
reg soc_videooverlaysoc_hdmi_in0_wer0_period_done = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer0_wer_counter = 24'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_r = 24'd0;
reg soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_r_updated = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_sys = 24'd0;
wire soc_videooverlaysoc_hdmi_in0_wer0_i;
wire soc_videooverlaysoc_hdmi_in0_wer0_o;
reg soc_videooverlaysoc_hdmi_in0_wer0_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_wer0_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_wer0_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_decoding0_valid_i;
wire [9:0] soc_videooverlaysoc_hdmi_in0_decoding0_input;
reg soc_videooverlaysoc_hdmi_in0_decoding0_valid_o = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in0_decoding0_output_raw = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_decoding0_output_d = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in0_decoding0_output_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in0_decoding0_output_de = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_d;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_re;
wire [4:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_r;
reg [4:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_w = 5'd0;
wire [1:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_status;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_phase_reset_re;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_phase_reset_r;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_phase_reset_w = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_i_nodelay;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_i_nodelay;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_rst;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_master_inc;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_master_ce;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_slave_inc;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_slave_ce;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_q;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_d;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_q;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_d;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
reg [9:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_o = 10'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst_write = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst_read = 1'd0;
wire hdmi_in0_data1_cap_write_clk;
wire hdmi_in0_data1_cap_write_rst;
wire hdmi_in0_data1_cap_read_clk;
wire hdmi_in0_data1_cap_read_rst;
reg [79:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr = 80'd0;
reg [79:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_rd = 80'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_wrpointer = 4'd5;
reg [2:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rdpointer = 3'd0;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_mdata;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_sdata;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_inc;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_dec;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_transition;
reg [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_mdata_d = 8'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture1_lateness = 8'd128;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_too_late;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_too_early;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_reset_lateness;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_charsync1_raw_data;
reg soc_videooverlaysoc_hdmi_in0_charsync1_synced = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in0_charsync1_data = 10'd0;
wire soc_videooverlaysoc_hdmi_in0_charsync1_char_synced_status;
wire [3:0] soc_videooverlaysoc_hdmi_in0_charsync1_ctl_pos_status;
reg [9:0] soc_videooverlaysoc_hdmi_in0_charsync1_raw_data1 = 10'd0;
wire [19:0] soc_videooverlaysoc_hdmi_in0_charsync1_raw;
reg soc_videooverlaysoc_hdmi_in0_charsync1_found_control = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_charsync1_control_position = 4'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in0_charsync1_control_counter = 3'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_charsync1_previous_control_position = 4'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_charsync1_word_sel = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_wer1_data;
wire soc_videooverlaysoc_hdmi_in0_wer1_update_re;
wire soc_videooverlaysoc_hdmi_in0_wer1_update_r;
reg soc_videooverlaysoc_hdmi_in0_wer1_update_w = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer1_status = 24'd0;
reg [8:0] soc_videooverlaysoc_hdmi_in0_wer1_data_r = 9'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_wer1_transitions = 8'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_wer1_transition_count = 4'd0;
reg soc_videooverlaysoc_hdmi_in0_wer1_is_control = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_wer1_is_error = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer1_period_counter = 24'd0;
reg soc_videooverlaysoc_hdmi_in0_wer1_period_done = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer1_wer_counter = 24'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_r = 24'd0;
reg soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_r_updated = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_sys = 24'd0;
wire soc_videooverlaysoc_hdmi_in0_wer1_i;
wire soc_videooverlaysoc_hdmi_in0_wer1_o;
reg soc_videooverlaysoc_hdmi_in0_wer1_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_wer1_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_wer1_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_decoding1_valid_i;
wire [9:0] soc_videooverlaysoc_hdmi_in0_decoding1_input;
reg soc_videooverlaysoc_hdmi_in0_decoding1_valid_o = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in0_decoding1_output_raw = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_decoding1_output_d = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in0_decoding1_output_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in0_decoding1_output_de = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_d;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_re;
wire [4:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_r;
reg [4:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_w = 5'd0;
wire [1:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_status;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_phase_reset_re;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_phase_reset_r;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_phase_reset_w = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_i_nodelay;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_i_nodelay;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_rst;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_master_inc;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_master_ce;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_slave_inc;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_slave_ce;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_q;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_d;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_q;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_d;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
reg [9:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_o = 10'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst_write = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst_read = 1'd0;
wire hdmi_in0_data2_cap_write_clk;
wire hdmi_in0_data2_cap_write_rst;
wire hdmi_in0_data2_cap_read_clk;
wire hdmi_in0_data2_cap_read_rst;
reg [79:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr = 80'd0;
reg [79:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_rd = 80'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_wrpointer = 4'd5;
reg [2:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rdpointer = 3'd0;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_mdata;
wire [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_sdata;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_inc;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_dec;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_transition;
reg [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_mdata_d = 8'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_s7datacapture2_lateness = 8'd128;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_too_late;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_too_early;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_reset_lateness;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_i;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_charsync2_raw_data;
reg soc_videooverlaysoc_hdmi_in0_charsync2_synced = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in0_charsync2_data = 10'd0;
wire soc_videooverlaysoc_hdmi_in0_charsync2_char_synced_status;
wire [3:0] soc_videooverlaysoc_hdmi_in0_charsync2_ctl_pos_status;
reg [9:0] soc_videooverlaysoc_hdmi_in0_charsync2_raw_data1 = 10'd0;
wire [19:0] soc_videooverlaysoc_hdmi_in0_charsync2_raw;
reg soc_videooverlaysoc_hdmi_in0_charsync2_found_control = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_charsync2_control_position = 4'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in0_charsync2_control_counter = 3'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_charsync2_previous_control_position = 4'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_charsync2_word_sel = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_wer2_data;
wire soc_videooverlaysoc_hdmi_in0_wer2_update_re;
wire soc_videooverlaysoc_hdmi_in0_wer2_update_r;
reg soc_videooverlaysoc_hdmi_in0_wer2_update_w = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer2_status = 24'd0;
reg [8:0] soc_videooverlaysoc_hdmi_in0_wer2_data_r = 9'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_wer2_transitions = 8'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_wer2_transition_count = 4'd0;
reg soc_videooverlaysoc_hdmi_in0_wer2_is_control = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_wer2_is_error = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer2_period_counter = 24'd0;
reg soc_videooverlaysoc_hdmi_in0_wer2_period_done = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer2_wer_counter = 24'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_r = 24'd0;
reg soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_r_updated = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_sys = 24'd0;
wire soc_videooverlaysoc_hdmi_in0_wer2_i;
wire soc_videooverlaysoc_hdmi_in0_wer2_o;
reg soc_videooverlaysoc_hdmi_in0_wer2_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_wer2_toggle_o;
reg soc_videooverlaysoc_hdmi_in0_wer2_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_decoding2_valid_i;
wire [9:0] soc_videooverlaysoc_hdmi_in0_decoding2_input;
reg soc_videooverlaysoc_hdmi_in0_decoding2_valid_o = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in0_decoding2_output_raw = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_decoding2_output_d = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in0_decoding2_output_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in0_decoding2_output_de = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_chansync_valid_i;
reg soc_videooverlaysoc_hdmi_in0_chansync_chan_synced = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_chansync_status;
wire soc_videooverlaysoc_hdmi_in0_chansync_all_control;
wire [9:0] soc_videooverlaysoc_hdmi_in0_chansync_data_in0_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_chansync_data_in0_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_chansync_data_in0_c;
wire soc_videooverlaysoc_hdmi_in0_chansync_data_in0_de;
wire [9:0] soc_videooverlaysoc_hdmi_in0_chansync_data_out0_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_chansync_data_out0_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_chansync_data_out0_c;
wire soc_videooverlaysoc_hdmi_in0_chansync_data_out0_de;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_din;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_dout;
wire soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_re;
reg [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_consume = 3'd0;
wire [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_dat_r;
wire soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_we;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_dat_w;
wire [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_rdport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_rdport_dat_r;
wire soc_videooverlaysoc_hdmi_in0_chansync_is_control0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_chansync_data_in1_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_chansync_data_in1_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_chansync_data_in1_c;
wire soc_videooverlaysoc_hdmi_in0_chansync_data_in1_de;
wire [9:0] soc_videooverlaysoc_hdmi_in0_chansync_data_out1_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_chansync_data_out1_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_chansync_data_out1_c;
wire soc_videooverlaysoc_hdmi_in0_chansync_data_out1_de;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_din;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_dout;
wire soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_re;
reg [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_consume = 3'd0;
wire [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_dat_r;
wire soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_we;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_dat_w;
wire [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_rdport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_rdport_dat_r;
wire soc_videooverlaysoc_hdmi_in0_chansync_is_control1;
wire [9:0] soc_videooverlaysoc_hdmi_in0_chansync_data_in2_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_chansync_data_in2_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_chansync_data_in2_c;
wire soc_videooverlaysoc_hdmi_in0_chansync_data_in2_de;
wire [9:0] soc_videooverlaysoc_hdmi_in0_chansync_data_out2_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_chansync_data_out2_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_chansync_data_out2_c;
wire soc_videooverlaysoc_hdmi_in0_chansync_data_out2_de;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_din;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_dout;
wire soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_re;
reg [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_consume = 3'd0;
wire [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_dat_r;
wire soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_we;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_dat_w;
wire [2:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_rdport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_rdport_dat_r;
wire soc_videooverlaysoc_hdmi_in0_chansync_is_control2;
wire soc_videooverlaysoc_hdmi_in0_chansync_some_control;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_valid_i;
wire [9:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_c;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_de;
wire [9:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_c;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_de;
wire [9:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_c;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_de;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_de_o = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_encoding_terc4 = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_storage_full = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_storage;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_dvimode_bit;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_de_r = 1'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_de = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_dgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_c;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_de;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_valid_in;
reg [1:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_de = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_c;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_de;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_valid_in;
reg [1:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_de = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_c;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_de;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_valid_in;
wire [3:0] soc_videooverlaysoc_hdmi_in0_decode_terc4_ctl_code;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_all_vgb;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_any_cvalid;
wire soc_videooverlaysoc_hdmi_in0_decode_terc4_c2c1_dgb;
wire soc_videooverlaysoc_hdmi_in0_syncpol_valid_i;
wire [9:0] soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_c;
wire soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_de;
wire [9:0] soc_videooverlaysoc_hdmi_in0_syncpol_data_in1_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_syncpol_data_in1_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_syncpol_data_in1_c;
wire soc_videooverlaysoc_hdmi_in0_syncpol_data_in1_de;
wire [9:0] soc_videooverlaysoc_hdmi_in0_syncpol_data_in2_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_syncpol_data_in2_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_syncpol_data_in2_c;
wire soc_videooverlaysoc_hdmi_in0_syncpol_data_in2_de;
reg soc_videooverlaysoc_hdmi_in0_syncpol_valid_o = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_syncpol_de;
wire soc_videooverlaysoc_hdmi_in0_syncpol_hsync;
wire soc_videooverlaysoc_hdmi_in0_syncpol_vsync;
reg [7:0] soc_videooverlaysoc_hdmi_in0_syncpol_r = 8'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_syncpol_g = 8'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_syncpol_b = 8'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in0_syncpol_c0 = 10'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in0_syncpol_c1 = 10'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in0_syncpol_c2 = 10'd0;
wire soc_videooverlaysoc_hdmi_in0_syncpol_de_rising;
wire soc_videooverlaysoc_hdmi_in0_syncpol_de_int;
reg soc_videooverlaysoc_hdmi_in0_syncpol_de_r = 1'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in0_syncpol_c_polarity = 2'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in0_syncpol_c_out = 2'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_c;
wire soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_de;
wire [9:0] soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_c;
wire soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_de;
reg [9:0] soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s0 = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s1 = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s2 = 2'd0;
reg soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s3 = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_c;
wire soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_de;
wire [9:0] soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_c;
wire soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_de;
reg [9:0] soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s0 = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s1 = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s2 = 2'd0;
reg soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s3 = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_c;
wire soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_de;
wire [9:0] soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_d;
wire [1:0] soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_c;
wire soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_de;
reg [9:0] soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s0 = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s1 = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s2 = 2'd0;
reg soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s3 = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_resdetection_valid_i;
wire soc_videooverlaysoc_hdmi_in0_resdetection_vsync;
wire soc_videooverlaysoc_hdmi_in0_resdetection_de;
wire [10:0] soc_videooverlaysoc_hdmi_in0_resdetection_hres_status;
wire [10:0] soc_videooverlaysoc_hdmi_in0_resdetection_vres_status;
reg soc_videooverlaysoc_hdmi_in0_resdetection_de_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_resdetection_pn_de;
reg [10:0] soc_videooverlaysoc_hdmi_in0_resdetection_hcounter = 11'd0;
reg [10:0] soc_videooverlaysoc_hdmi_in0_resdetection_hcounter_st = 11'd0;
reg soc_videooverlaysoc_hdmi_in0_resdetection_vsync_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_resdetection_p_vsync;
reg [10:0] soc_videooverlaysoc_hdmi_in0_resdetection_vcounter = 11'd0;
reg [10:0] soc_videooverlaysoc_hdmi_in0_resdetection_vcounter_st = 11'd0;
wire [9:0] soc_videooverlaysoc_hdmi_out0_clk_gen_data0;
wire [9:0] soc_videooverlaysoc_hdmi_out0_clk_gen_data1;
reg soc_videooverlaysoc_hdmi_out0_clk_gen_ce = 1'd0;
wire [1:0] soc_videooverlaysoc_hdmi_out0_clk_gen_shift;
wire soc_videooverlaysoc_hdmi_out0_clk_gen_pad_se;
reg [9:0] soc_videooverlaysoc = 10'd31;
wire soc_videooverlaysoc_hdmi_out0_phy_sink_ready;
reg [9:0] soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c0 = 10'd0;
reg [9:0] soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c1 = 10'd0;
reg [10:0] soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c2 = 11'd0;
wire [9:0] soc_videooverlaysoc_hdmi_out0_phy_es0_data0;
wire [9:0] soc_videooverlaysoc_hdmi_out0_phy_es0_data1;
reg soc_videooverlaysoc_hdmi_out0_phy_es0_ce = 1'd0;
wire [1:0] soc_videooverlaysoc_hdmi_out0_phy_es0_shift;
wire soc_videooverlaysoc_hdmi_out0_phy_es0_pad_se;
wire [9:0] soc_videooverlaysoc_hdmi_out0_phy_es1_data0;
wire [9:0] soc_videooverlaysoc_hdmi_out0_phy_es1_data1;
reg soc_videooverlaysoc_hdmi_out0_phy_es1_ce = 1'd0;
wire [1:0] soc_videooverlaysoc_hdmi_out0_phy_es1_shift;
wire soc_videooverlaysoc_hdmi_out0_phy_es1_pad_se;
wire [9:0] soc_videooverlaysoc_hdmi_out0_phy_es2_data0;
wire [9:0] soc_videooverlaysoc_hdmi_out0_phy_es2_data1;
reg soc_videooverlaysoc_hdmi_out0_phy_es2_ce = 1'd0;
wire [1:0] soc_videooverlaysoc_hdmi_out0_phy_es2_shift;
wire soc_videooverlaysoc_hdmi_out0_phy_es2_pad_se;
reg soc_videooverlaysoc_hdmi_in0_timing_valid = 1'd0;
wire soc_videooverlaysoc_hdmi_in0_timing_ready;
reg soc_videooverlaysoc_hdmi_in0_timing_first = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_timing_last = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_timing_payload_hsync = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_timing_payload_vsync = 1'd0;
reg soc_videooverlaysoc_hdmi_in0_timing_payload_de = 1'd0;
wire soc_videooverlaysoc_early_line_end;
wire soc_videooverlaysoc_hdmi_in1_freq_clk0;
wire [31:0] soc_videooverlaysoc_hdmi_in1_freq_status;
wire hdmi_in1_freq_fmeter_clk;
wire soc_videooverlaysoc_hdmi_in1_freq_period_done;
reg [31:0] soc_videooverlaysoc_hdmi_in1_freq_period_counter = 32'd0;
wire soc_videooverlaysoc_hdmi_in1_freq_ce;
reg [5:0] soc_videooverlaysoc_hdmi_in1_freq_q = 6'd0;
wire [5:0] soc_videooverlaysoc_hdmi_in1_freq_q_next;
reg [5:0] soc_videooverlaysoc_hdmi_in1_freq_q_binary = 6'd0;
reg [5:0] soc_videooverlaysoc_hdmi_in1_freq_q_next_binary = 6'd0;
wire [5:0] soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_i;
reg [5:0] soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o = 6'd0;
reg [5:0] soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb = 6'd0;
wire soc_videooverlaysoc_hdmi_in1_freq_sampler_latch;
wire [5:0] soc_videooverlaysoc_hdmi_in1_freq_sampler_i;
reg [31:0] soc_videooverlaysoc_hdmi_in1_freq_sampler_o = 32'd0;
wire [5:0] soc_videooverlaysoc_hdmi_in1_freq_sampler_inc;
reg [31:0] soc_videooverlaysoc_hdmi_in1_freq_sampler_counter = 32'd0;
reg [5:0] soc_videooverlaysoc_hdmi_in1_freq_sampler_i_d = 6'd0;
wire soc_videooverlaysoc_litedramcrossbar_cmd_valid;
wire soc_videooverlaysoc_litedramcrossbar_cmd_ready;
wire soc_videooverlaysoc_litedramcrossbar_cmd_payload_we;
wire [23:0] soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr;
wire soc_videooverlaysoc_litedramcrossbar_wdata_valid;
wire soc_videooverlaysoc_litedramcrossbar_wdata_ready;
wire [255:0] soc_videooverlaysoc_litedramcrossbar_wdata_payload_data;
wire [31:0] soc_videooverlaysoc_litedramcrossbar_wdata_payload_we;
wire soc_videooverlaysoc_litedramcrossbar_rdata_valid;
wire [255:0] soc_videooverlaysoc_litedramcrossbar_rdata_payload_data;
wire soc_videooverlaysoc_hdmi_in1_edid_status;
reg soc_videooverlaysoc_hdmi_in1_edid_storage_full = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_edid_storage;
reg soc_videooverlaysoc_hdmi_in1_edid_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_edid_scl_raw;
reg soc_videooverlaysoc_hdmi_in1_edid_sda_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_edid_sda_raw;
reg soc_videooverlaysoc_hdmi_in1_edid_sda_drv = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_sda_drv_reg = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_edid_sda_i_async;
wire soc_videooverlaysoc_hdmi_in1_edid_sda_o;
reg soc_videooverlaysoc_hdmi_in1_edid_scl_i = 1'd0;
reg [5:0] soc_videooverlaysoc_hdmi_in1_edid_samp_count = 6'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_samp_carry = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_scl_r = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_sda_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_edid_scl_rising;
wire soc_videooverlaysoc_hdmi_in1_edid_sda_rising;
wire soc_videooverlaysoc_hdmi_in1_edid_sda_falling;
wire soc_videooverlaysoc_hdmi_in1_edid_start;
reg [7:0] soc_videooverlaysoc_hdmi_in1_edid_din = 8'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_edid_counter = 4'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_is_read = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_update_is_read = 1'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_edid_offset_counter = 8'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_oc_load = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_oc_inc = 1'd0;
wire [7:0] soc_videooverlaysoc_hdmi_in1_edid_adr;
wire [7:0] soc_videooverlaysoc_hdmi_in1_edid_dat_r;
reg soc_videooverlaysoc_hdmi_in1_edid_data_bit = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_zero_drv = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_data_drv = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_data_drv_en = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_edid_data_drv_stop = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_mmcm_reset_storage_full = 1'd1;
wire soc_videooverlaysoc_hdmi_in1_mmcm_reset_storage;
reg soc_videooverlaysoc_hdmi_in1_mmcm_reset_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_locked_status;
wire soc_videooverlaysoc_hdmi_in1_mmcm_read_re;
wire soc_videooverlaysoc_hdmi_in1_mmcm_read_r;
reg soc_videooverlaysoc_hdmi_in1_mmcm_read_w = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_mmcm_write_re;
wire soc_videooverlaysoc_hdmi_in1_mmcm_write_r;
reg soc_videooverlaysoc_hdmi_in1_mmcm_write_w = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_mmcm_drdy_status = 1'd0;
reg [6:0] soc_videooverlaysoc_hdmi_in1_mmcm_adr_storage_full = 7'd0;
wire [6:0] soc_videooverlaysoc_hdmi_in1_mmcm_adr_storage;
reg soc_videooverlaysoc_hdmi_in1_mmcm_adr_re = 1'd0;
reg [15:0] soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_storage_full = 16'd0;
wire [15:0] soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_storage;
reg soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_re = 1'd0;
wire [15:0] soc_videooverlaysoc_hdmi_in1_mmcm_dat_r_status;
wire soc_videooverlaysoc_hdmi_in1_locked;
wire hdmi_in1_pix_clk;
wire hdmi_in1_pix_rst;
wire hdmi_in1_pix1p25x_clk;
wire hdmi_in1_pix1p25x_rst;
wire hdmi_in1_pix5x_clk;
wire soc_videooverlaysoc_hdmi_in1_clk_input;
wire soc_videooverlaysoc_hdmi_in1_clk_input_bufr;
wire soc_videooverlaysoc_hdmi_in1_mmcm_fb;
wire soc_videooverlaysoc_hdmi_in1_mmcm_locked;
wire soc_videooverlaysoc_hdmi_in1_mmcm_clk0;
wire soc_videooverlaysoc_hdmi_in1_mmcm_clk1;
wire soc_videooverlaysoc_hdmi_in1_mmcm_clk2;
wire soc_videooverlaysoc_hdmi_in1_mmcm_drdy;
wire soc_videooverlaysoc_hdmi_in1_mmcm_fb_o;
wire [9:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_d;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_re;
wire [4:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_r;
reg [4:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_w = 5'd0;
wire [1:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_status;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_phase_reset_re;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_phase_reset_r;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_phase_reset_w = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_i_nodelay;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_i_nodelay;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_rst;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_master_inc;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_master_ce;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_slave_inc;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_slave_ce;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_q;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_d;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_q;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_d;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
reg [9:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_o = 10'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst_write = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst_read = 1'd0;
wire hdmi_in1_data0_cap_write_clk;
wire hdmi_in1_data0_cap_write_rst;
wire hdmi_in1_data0_cap_read_clk;
wire hdmi_in1_data0_cap_read_rst;
reg [79:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr = 80'd0;
reg [79:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_rd = 80'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_wrpointer = 4'd5;
reg [2:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rdpointer = 3'd0;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_mdata;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_sdata;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_inc;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_dec;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_transition;
reg [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_mdata_d = 8'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture0_lateness = 8'd128;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_too_late;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_too_early;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_reset_lateness;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_charsync0_raw_data;
reg soc_videooverlaysoc_hdmi_in1_charsync0_synced = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in1_charsync0_data = 10'd0;
wire soc_videooverlaysoc_hdmi_in1_charsync0_char_synced_status;
wire [3:0] soc_videooverlaysoc_hdmi_in1_charsync0_ctl_pos_status;
reg [9:0] soc_videooverlaysoc_hdmi_in1_charsync0_raw_data1 = 10'd0;
wire [19:0] soc_videooverlaysoc_hdmi_in1_charsync0_raw;
reg soc_videooverlaysoc_hdmi_in1_charsync0_found_control = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_charsync0_control_position = 4'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in1_charsync0_control_counter = 3'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_charsync0_previous_control_position = 4'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_charsync0_word_sel = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_wer0_data;
wire soc_videooverlaysoc_hdmi_in1_wer0_update_re;
wire soc_videooverlaysoc_hdmi_in1_wer0_update_r;
reg soc_videooverlaysoc_hdmi_in1_wer0_update_w = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer0_status = 24'd0;
reg [8:0] soc_videooverlaysoc_hdmi_in1_wer0_data_r = 9'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_wer0_transitions = 8'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_wer0_transition_count = 4'd0;
reg soc_videooverlaysoc_hdmi_in1_wer0_is_control = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_wer0_is_error = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer0_period_counter = 24'd0;
reg soc_videooverlaysoc_hdmi_in1_wer0_period_done = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer0_wer_counter = 24'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_r = 24'd0;
reg soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_r_updated = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_sys = 24'd0;
wire soc_videooverlaysoc_hdmi_in1_wer0_i;
wire soc_videooverlaysoc_hdmi_in1_wer0_o;
reg soc_videooverlaysoc_hdmi_in1_wer0_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_wer0_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_wer0_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_decoding0_valid_i;
wire [9:0] soc_videooverlaysoc_hdmi_in1_decoding0_input;
reg soc_videooverlaysoc_hdmi_in1_decoding0_valid_o = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in1_decoding0_output_raw = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_decoding0_output_d = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in1_decoding0_output_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in1_decoding0_output_de = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_d;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_re;
wire [4:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_r;
reg [4:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_w = 5'd0;
wire [1:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_status;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_phase_reset_re;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_phase_reset_r;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_phase_reset_w = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_i_nodelay;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_i_nodelay;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_rst;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_master_inc;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_master_ce;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_slave_inc;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_slave_ce;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_q;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_d;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_q;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_d;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
reg [9:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_o = 10'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst_write = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst_read = 1'd0;
wire hdmi_in1_data1_cap_write_clk;
wire hdmi_in1_data1_cap_write_rst;
wire hdmi_in1_data1_cap_read_clk;
wire hdmi_in1_data1_cap_read_rst;
reg [79:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr = 80'd0;
reg [79:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_rd = 80'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_wrpointer = 4'd5;
reg [2:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rdpointer = 3'd0;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_mdata;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_sdata;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_inc;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_dec;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_transition;
reg [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_mdata_d = 8'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture1_lateness = 8'd128;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_too_late;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_too_early;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_reset_lateness;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_charsync1_raw_data;
reg soc_videooverlaysoc_hdmi_in1_charsync1_synced = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in1_charsync1_data = 10'd0;
wire soc_videooverlaysoc_hdmi_in1_charsync1_char_synced_status;
wire [3:0] soc_videooverlaysoc_hdmi_in1_charsync1_ctl_pos_status;
reg [9:0] soc_videooverlaysoc_hdmi_in1_charsync1_raw_data1 = 10'd0;
wire [19:0] soc_videooverlaysoc_hdmi_in1_charsync1_raw;
reg soc_videooverlaysoc_hdmi_in1_charsync1_found_control = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_charsync1_control_position = 4'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in1_charsync1_control_counter = 3'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_charsync1_previous_control_position = 4'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_charsync1_word_sel = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_wer1_data;
wire soc_videooverlaysoc_hdmi_in1_wer1_update_re;
wire soc_videooverlaysoc_hdmi_in1_wer1_update_r;
reg soc_videooverlaysoc_hdmi_in1_wer1_update_w = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer1_status = 24'd0;
reg [8:0] soc_videooverlaysoc_hdmi_in1_wer1_data_r = 9'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_wer1_transitions = 8'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_wer1_transition_count = 4'd0;
reg soc_videooverlaysoc_hdmi_in1_wer1_is_control = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_wer1_is_error = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer1_period_counter = 24'd0;
reg soc_videooverlaysoc_hdmi_in1_wer1_period_done = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer1_wer_counter = 24'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_r = 24'd0;
reg soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_r_updated = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_sys = 24'd0;
wire soc_videooverlaysoc_hdmi_in1_wer1_i;
wire soc_videooverlaysoc_hdmi_in1_wer1_o;
reg soc_videooverlaysoc_hdmi_in1_wer1_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_wer1_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_wer1_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_decoding1_valid_i;
wire [9:0] soc_videooverlaysoc_hdmi_in1_decoding1_input;
reg soc_videooverlaysoc_hdmi_in1_decoding1_valid_o = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in1_decoding1_output_raw = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_decoding1_output_d = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in1_decoding1_output_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in1_decoding1_output_de = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_d;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_re;
wire [4:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_r;
reg [4:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_w = 5'd0;
wire [1:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_status;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_phase_reset_re;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_phase_reset_r;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_phase_reset_w = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_i_nodelay;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_i_nodelay;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_rst;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_master_inc;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_master_ce;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_slave_inc;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_slave_ce;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_q;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_d;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_i_delayed;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_q;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_d;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
reg [9:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_o = 10'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst_write = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst_read = 1'd0;
wire hdmi_in1_data2_cap_write_clk;
wire hdmi_in1_data2_cap_write_rst;
wire hdmi_in1_data2_cap_read_clk;
wire hdmi_in1_data2_cap_read_rst;
reg [79:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr = 80'd0;
reg [79:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_rd = 80'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_wrpointer = 4'd5;
reg [2:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rdpointer = 3'd0;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_mdata;
wire [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_sdata;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_inc;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_dec;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_transition;
reg [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_mdata_d = 8'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_s7datacapture2_lateness = 8'd128;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_too_late;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_too_early;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_reset_lateness;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_i;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_charsync2_raw_data;
reg soc_videooverlaysoc_hdmi_in1_charsync2_synced = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in1_charsync2_data = 10'd0;
wire soc_videooverlaysoc_hdmi_in1_charsync2_char_synced_status;
wire [3:0] soc_videooverlaysoc_hdmi_in1_charsync2_ctl_pos_status;
reg [9:0] soc_videooverlaysoc_hdmi_in1_charsync2_raw_data1 = 10'd0;
wire [19:0] soc_videooverlaysoc_hdmi_in1_charsync2_raw;
reg soc_videooverlaysoc_hdmi_in1_charsync2_found_control = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_charsync2_control_position = 4'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in1_charsync2_control_counter = 3'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_charsync2_previous_control_position = 4'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_charsync2_word_sel = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_wer2_data;
wire soc_videooverlaysoc_hdmi_in1_wer2_update_re;
wire soc_videooverlaysoc_hdmi_in1_wer2_update_r;
reg soc_videooverlaysoc_hdmi_in1_wer2_update_w = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer2_status = 24'd0;
reg [8:0] soc_videooverlaysoc_hdmi_in1_wer2_data_r = 9'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_wer2_transitions = 8'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_wer2_transition_count = 4'd0;
reg soc_videooverlaysoc_hdmi_in1_wer2_is_control = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_wer2_is_error = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer2_period_counter = 24'd0;
reg soc_videooverlaysoc_hdmi_in1_wer2_period_done = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer2_wer_counter = 24'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_r = 24'd0;
reg soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_r_updated = 1'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_sys = 24'd0;
wire soc_videooverlaysoc_hdmi_in1_wer2_i;
wire soc_videooverlaysoc_hdmi_in1_wer2_o;
reg soc_videooverlaysoc_hdmi_in1_wer2_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_wer2_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_wer2_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_decoding2_valid_i;
wire [9:0] soc_videooverlaysoc_hdmi_in1_decoding2_input;
reg soc_videooverlaysoc_hdmi_in1_decoding2_valid_o = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in1_decoding2_output_raw = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_decoding2_output_d = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in1_decoding2_output_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in1_decoding2_output_de = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_chansync_valid_i;
reg soc_videooverlaysoc_hdmi_in1_chansync_chan_synced = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_chansync_status;
wire soc_videooverlaysoc_hdmi_in1_chansync_all_control;
wire [9:0] soc_videooverlaysoc_hdmi_in1_chansync_data_in0_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_chansync_data_in0_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_chansync_data_in0_c;
wire soc_videooverlaysoc_hdmi_in1_chansync_data_in0_de;
wire [9:0] soc_videooverlaysoc_hdmi_in1_chansync_data_out0_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_chansync_data_out0_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_chansync_data_out0_c;
wire soc_videooverlaysoc_hdmi_in1_chansync_data_out0_de;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_din;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_dout;
wire soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_re;
reg [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_consume = 3'd0;
wire [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_dat_r;
wire soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_we;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_dat_w;
wire [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_rdport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_rdport_dat_r;
wire soc_videooverlaysoc_hdmi_in1_chansync_is_control0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_chansync_data_in1_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_chansync_data_in1_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_chansync_data_in1_c;
wire soc_videooverlaysoc_hdmi_in1_chansync_data_in1_de;
wire [9:0] soc_videooverlaysoc_hdmi_in1_chansync_data_out1_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_chansync_data_out1_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_chansync_data_out1_c;
wire soc_videooverlaysoc_hdmi_in1_chansync_data_out1_de;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_din;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_dout;
wire soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_re;
reg [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_consume = 3'd0;
wire [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_dat_r;
wire soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_we;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_dat_w;
wire [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_rdport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_rdport_dat_r;
wire soc_videooverlaysoc_hdmi_in1_chansync_is_control1;
wire [9:0] soc_videooverlaysoc_hdmi_in1_chansync_data_in2_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_chansync_data_in2_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_chansync_data_in2_c;
wire soc_videooverlaysoc_hdmi_in1_chansync_data_in2_de;
wire [9:0] soc_videooverlaysoc_hdmi_in1_chansync_data_out2_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_chansync_data_out2_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_chansync_data_out2_c;
wire soc_videooverlaysoc_hdmi_in1_chansync_data_out2_de;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_din;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_dout;
wire soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_re;
reg [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_consume = 3'd0;
wire [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_dat_r;
wire soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_we;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_dat_w;
wire [2:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_rdport_adr;
wire [20:0] soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_rdport_dat_r;
wire soc_videooverlaysoc_hdmi_in1_chansync_is_control2;
wire soc_videooverlaysoc_hdmi_in1_chansync_some_control;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_valid_i;
wire [9:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_c;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_de;
wire [9:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_c;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_de;
wire [9:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_c;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_de;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_de_o = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_encoding_terc4 = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_video = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_data = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_storage_full = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_storage;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_dvimode_bit;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_de_r = 1'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_de = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_dgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_c;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_de;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_valid_in;
reg [1:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_de = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_c;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_de;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_valid_in;
reg [1:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c = 2'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_de = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d = 4'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_c;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_de;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_valid_in;
wire [3:0] soc_videooverlaysoc_hdmi_in1_decode_terc4_ctl_code;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_all_vgb;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_any_cvalid;
wire soc_videooverlaysoc_hdmi_in1_decode_terc4_c2c1_dgb;
wire soc_videooverlaysoc_hdmi_in1_syncpol_valid_i;
wire [9:0] soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_c;
wire soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_de;
wire [9:0] soc_videooverlaysoc_hdmi_in1_syncpol_data_in1_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_syncpol_data_in1_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_syncpol_data_in1_c;
wire soc_videooverlaysoc_hdmi_in1_syncpol_data_in1_de;
wire [9:0] soc_videooverlaysoc_hdmi_in1_syncpol_data_in2_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_syncpol_data_in2_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_syncpol_data_in2_c;
wire soc_videooverlaysoc_hdmi_in1_syncpol_data_in2_de;
reg soc_videooverlaysoc_hdmi_in1_syncpol_valid_o = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_syncpol_de;
wire soc_videooverlaysoc_hdmi_in1_syncpol_hsync;
wire soc_videooverlaysoc_hdmi_in1_syncpol_vsync;
reg [7:0] soc_videooverlaysoc_hdmi_in1_syncpol_r = 8'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_syncpol_g = 8'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_syncpol_b = 8'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in1_syncpol_c0 = 10'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in1_syncpol_c1 = 10'd0;
reg [9:0] soc_videooverlaysoc_hdmi_in1_syncpol_c2 = 10'd0;
wire soc_videooverlaysoc_hdmi_in1_syncpol_de_rising;
wire soc_videooverlaysoc_hdmi_in1_syncpol_de_int;
reg soc_videooverlaysoc_hdmi_in1_syncpol_de_r = 1'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in1_syncpol_c_polarity = 2'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in1_syncpol_c_out = 2'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_c;
wire soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_de;
wire [9:0] soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_c;
wire soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_de;
reg [9:0] soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s0 = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s1 = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s2 = 2'd0;
reg soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s3 = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_c;
wire soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_de;
wire [9:0] soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_c;
wire soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_de;
reg [9:0] soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s0 = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s1 = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s2 = 2'd0;
reg soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s3 = 1'd0;
wire [9:0] soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_c;
wire soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_de;
wire [9:0] soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_raw;
wire [7:0] soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_d;
wire [1:0] soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_c;
wire soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_de;
reg [9:0] soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s0 = 10'd0;
reg [7:0] soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s1 = 8'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s2 = 2'd0;
reg soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s3 = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_resdetection_valid_i;
wire soc_videooverlaysoc_hdmi_in1_resdetection_vsync;
wire soc_videooverlaysoc_hdmi_in1_resdetection_de;
wire [10:0] soc_videooverlaysoc_hdmi_in1_resdetection_hres_status;
wire [10:0] soc_videooverlaysoc_hdmi_in1_resdetection_vres_status;
reg soc_videooverlaysoc_hdmi_in1_resdetection_de_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_resdetection_pn_de;
reg [10:0] soc_videooverlaysoc_hdmi_in1_resdetection_hcounter = 11'd0;
reg [10:0] soc_videooverlaysoc_hdmi_in1_resdetection_hcounter_st = 11'd0;
reg soc_videooverlaysoc_hdmi_in1_resdetection_vsync_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_resdetection_p_vsync;
reg [10:0] soc_videooverlaysoc_hdmi_in1_resdetection_vcounter = 11'd0;
reg [10:0] soc_videooverlaysoc_hdmi_in1_resdetection_vcounter_st = 11'd0;
wire soc_videooverlaysoc_hdmi_in1_frame_valid_i;
wire soc_videooverlaysoc_hdmi_in1_frame_vsync;
wire soc_videooverlaysoc_hdmi_in1_frame_de;
wire [7:0] soc_videooverlaysoc_hdmi_in1_frame_r;
wire [7:0] soc_videooverlaysoc_hdmi_in1_frame_g;
wire [7:0] soc_videooverlaysoc_hdmi_in1_frame_b;
wire soc_videooverlaysoc_hdmi_in1_frame_frame_valid;
wire soc_videooverlaysoc_hdmi_in1_frame_frame_ready;
wire soc_videooverlaysoc_hdmi_in1_frame_frame_first;
wire soc_videooverlaysoc_hdmi_in1_frame_frame_last;
wire soc_videooverlaysoc_hdmi_in1_frame_frame_payload_sof;
wire [255:0] soc_videooverlaysoc_hdmi_in1_frame_frame_payload_pixels;
wire soc_videooverlaysoc_hdmi_in1_frame_busy;
wire soc_videooverlaysoc_hdmi_in1_frame_overflow_re;
wire soc_videooverlaysoc_hdmi_in1_frame_overflow_r;
wire soc_videooverlaysoc_hdmi_in1_frame_overflow_w;
reg soc_videooverlaysoc_hdmi_in1_frame_vsync_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_frame_new_frame;
reg [255:0] soc_videooverlaysoc_hdmi_in1_frame_cur_word = 256'd0;
reg soc_videooverlaysoc_hdmi_in1_frame_cur_word_valid = 1'd0;
wire [31:0] soc_videooverlaysoc_hdmi_in1_frame_encoded_pixel;
reg [7:0] soc_videooverlaysoc_hdmi_in1_frame_dummy8 = 8'd0;
reg [2:0] soc_videooverlaysoc_hdmi_in1_frame_pack_counter = 3'd0;
wire soc_videooverlaysoc_hdmi_in1_frame_sink_valid;
wire soc_videooverlaysoc_hdmi_in1_frame_sink_ready;
reg soc_videooverlaysoc_hdmi_in1_frame_sink_first = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_frame_sink_last = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_frame_sink_payload_sof = 1'd0;
wire [255:0] soc_videooverlaysoc_hdmi_in1_frame_sink_payload_pixels;
wire soc_videooverlaysoc_hdmi_in1_frame_source_valid;
wire soc_videooverlaysoc_hdmi_in1_frame_source_ready;
wire soc_videooverlaysoc_hdmi_in1_frame_source_first;
wire soc_videooverlaysoc_hdmi_in1_frame_source_last;
wire soc_videooverlaysoc_hdmi_in1_frame_source_payload_sof;
wire [255:0] soc_videooverlaysoc_hdmi_in1_frame_source_payload_pixels;
wire soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_we;
wire soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_writable;
wire soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_re;
wire soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_readable;
wire [258:0] soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_din;
wire [258:0] soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_dout;
wire soc_videooverlaysoc_hdmi_in1_frame_graycounter0_ce;
(* dont_touch = "true" *) reg [10:0] soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q = 11'd0;
wire [10:0] soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_next;
reg [10:0] soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_binary = 11'd0;
reg [10:0] soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_next_binary = 11'd0;
wire soc_videooverlaysoc_hdmi_in1_frame_graycounter1_ce;
(* dont_touch = "true" *) reg [10:0] soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q = 11'd0;
wire [10:0] soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next;
reg [10:0] soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_binary = 11'd0;
reg [10:0] soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next_binary = 11'd0;
wire [10:0] soc_videooverlaysoc_hdmi_in1_frame_produce_rdomain;
wire [10:0] soc_videooverlaysoc_hdmi_in1_frame_consume_wdomain;
wire [9:0] soc_videooverlaysoc_hdmi_in1_frame_wrport_adr;
wire [258:0] soc_videooverlaysoc_hdmi_in1_frame_wrport_dat_r;
wire soc_videooverlaysoc_hdmi_in1_frame_wrport_we;
wire [258:0] soc_videooverlaysoc_hdmi_in1_frame_wrport_dat_w;
wire [9:0] soc_videooverlaysoc_hdmi_in1_frame_rdport_adr;
wire [258:0] soc_videooverlaysoc_hdmi_in1_frame_rdport_dat_r;
wire soc_videooverlaysoc_hdmi_in1_frame_fifo_in_payload_sof;
wire [255:0] soc_videooverlaysoc_hdmi_in1_frame_fifo_in_payload_pixels;
wire soc_videooverlaysoc_hdmi_in1_frame_fifo_in_first;
wire soc_videooverlaysoc_hdmi_in1_frame_fifo_in_last;
wire soc_videooverlaysoc_hdmi_in1_frame_fifo_out_payload_sof;
wire [255:0] soc_videooverlaysoc_hdmi_in1_frame_fifo_out_payload_pixels;
wire soc_videooverlaysoc_hdmi_in1_frame_fifo_out_first;
wire soc_videooverlaysoc_hdmi_in1_frame_fifo_out_last;
reg soc_videooverlaysoc_hdmi_in1_frame_pix_overflow = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_frame_pix_overflow_reset;
wire soc_videooverlaysoc_hdmi_in1_frame_sys_overflow;
wire soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_i;
wire soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_o;
reg soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_i;
wire soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_o;
reg soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_o;
reg soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_o_r = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_frame_overflow_mask = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_frame_valid;
reg soc_videooverlaysoc_hdmi_in1_dma_frame_ready = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_frame_first;
wire soc_videooverlaysoc_hdmi_in1_dma_frame_last;
wire soc_videooverlaysoc_hdmi_in1_dma_frame_payload_sof;
wire [255:0] soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels;
reg [28:0] soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full = 29'd0;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage;
reg soc_videooverlaysoc_hdmi_in1_dma_frame_size_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_irq;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_address;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_reached;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_valid;
reg soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_done = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_pending;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_trigger;
reg soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_clear = 1'd0;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_reached;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_valid;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_done;
reg [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_storage_full = 2'd0;
wire [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_storage;
reg soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_we;
wire [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_dat_w;
reg [28:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full = 29'd0;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage;
reg soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_we;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_dat_w;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_pending;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_trigger;
reg soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_clear = 1'd0;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_reached;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_valid;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_done;
reg [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_storage_full = 2'd0;
wire [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_storage;
reg soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_we;
wire [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_dat_w;
reg [28:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full = 29'd0;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage;
reg soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_we;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_dat_w;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_status_re;
wire [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_status_r;
reg [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_status_w = 2'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_re;
wire [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_r;
reg [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_w = 2'd0;
reg [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_storage_full = 2'd0;
wire [1:0] soc_videooverlaysoc_hdmi_in1_dma_slot_array_storage;
reg soc_videooverlaysoc_hdmi_in1_dma_slot_array_re = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_slot_array_change_slot;
reg soc_videooverlaysoc_hdmi_in1_dma_slot_array_current_slot = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_dma_reset_words = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_dma_count_word = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_last_word;
reg [23:0] soc_videooverlaysoc_hdmi_in1_dma_current_address = 24'd0;
reg [23:0] soc_videooverlaysoc_hdmi_in1_dma_mwords_remaining = 24'd0;
wire [255:0] soc_videooverlaysoc_hdmi_in1_dma_memory_word;
reg soc_videooverlaysoc_hdmi_in1_dma_sink_sink_valid = 1'd0;
wire soc_videooverlaysoc_hdmi_in1_dma_sink_sink_ready;
wire [23:0] soc_videooverlaysoc_hdmi_in1_dma_sink_sink_payload_address;
wire [255:0] soc_videooverlaysoc_hdmi_in1_dma_sink_sink_payload_data;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_valid;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_ready;
reg soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_first = 1'd0;
reg soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_last = 1'd0;
wire [255:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_payload_data;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_source_valid;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_source_ready;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_source_first;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_source_last;
wire [255:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_source_payload_data;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_we;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_writable;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_re;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_readable;
wire [257:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_din;
wire [257:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_dout;
reg [4:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_level = 5'd0;
reg soc_videooverlaysoc_hdmi_in1_dma_fifo_replace = 1'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_produce = 4'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_consume = 4'd0;
reg [3:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_adr = 4'd0;
wire [257:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_dat_r;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_we;
wire [257:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_dat_w;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_do_read;
wire [3:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_rdport_adr;
wire [257:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_rdport_dat_r;
wire [255:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_in_payload_data;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_in_first;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_in_last;
wire [255:0] soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_out_payload_data;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_out_first;
wire soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_out_last;
wire soc_videooverlaysoc_out_dram_port_cmd_valid;
wire soc_videooverlaysoc_out_dram_port_cmd_ready;
wire soc_videooverlaysoc_out_dram_port_cmd_first;
wire soc_videooverlaysoc_out_dram_port_cmd_last;
wire soc_videooverlaysoc_out_dram_port_cmd_payload_we;
wire [23:0] soc_videooverlaysoc_out_dram_port_cmd_payload_addr;
wire soc_videooverlaysoc_out_dram_port_wdata_ready;
reg [255:0] soc_videooverlaysoc_out_dram_port_wdata_payload_data = 256'd0;
reg [31:0] soc_videooverlaysoc_out_dram_port_wdata_payload_we = 32'd0;
wire soc_videooverlaysoc_out_dram_port_rdata_valid;
wire soc_videooverlaysoc_out_dram_port_rdata_ready;
reg soc_videooverlaysoc_out_dram_port_rdata_first = 1'd0;
reg soc_videooverlaysoc_out_dram_port_rdata_last = 1'd0;
wire [255:0] soc_videooverlaysoc_out_dram_port_rdata_payload_data;
reg soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_valid = 1'd0;
wire soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_ready;
reg soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_first = 1'd0;
reg soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_last = 1'd0;
reg soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_payload_we = 1'd0;
reg [23:0] soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_payload_addr = 24'd0;
wire soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_valid;
wire soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_ready;
wire soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_first;
wire soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_last;
wire [255:0] soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_payload_data;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_valid;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_ready;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_first;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_last;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_payload_we;
wire [23:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_payload_addr;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_source_valid;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_source_ready;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_source_first;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_source_last;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_source_payload_we;
wire [23:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_source_payload_addr;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_we;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_writable;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_re;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_readable;
wire [26:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_din;
wire [26:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_dout;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_ce;
(* dont_touch = "true" *) reg [2:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q = 3'd0;
wire [2:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_next;
reg [2:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_binary = 3'd0;
reg [2:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_next_binary = 3'd0;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_ce;
(* dont_touch = "true" *) reg [2:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q = 3'd0;
wire [2:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next;
reg [2:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_binary = 3'd0;
reg [2:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next_binary = 3'd0;
wire [2:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_produce_rdomain;
wire [2:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_consume_wdomain;
wire [1:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_adr;
wire [26:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_dat_r;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_we;
wire [26:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_dat_w;
wire [1:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_rdport_adr;
wire [26:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_rdport_dat_r;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_payload_we;
wire [23:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_payload_addr;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_first;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_last;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_payload_we;
wire [23:0] soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_payload_addr;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_first;
wire soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_last;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_valid;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_ready;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_first;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_last;
wire [255:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_payload_data;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_source_valid;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_source_ready;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_source_first;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_source_last;
wire [255:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_source_payload_data;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_we;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_writable;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_re;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_readable;
wire [257:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_din;
wire [257:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_dout;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_ce;
(* dont_touch = "true" *) reg [4:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q = 5'd0;
wire [4:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_next;
reg [4:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_binary = 5'd0;
reg [4:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_next_binary = 5'd0;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_ce;
(* dont_touch = "true" *) reg [4:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q = 5'd0;
wire [4:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next;
reg [4:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_binary = 5'd0;
reg [4:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next_binary = 5'd0;
wire [4:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_produce_rdomain;
wire [4:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_consume_wdomain;
wire [3:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_adr;
wire [257:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_dat_r;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_we;
wire [257:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_dat_w;
wire [3:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_rdport_adr;
wire [257:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_rdport_dat_r;
wire [255:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_in_payload_data;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_in_first;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_in_last;
wire [255:0] soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_out_payload_data;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_out_first;
wire soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_out_last;
wire soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_valid;
reg soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_ready = 1'd0;
wire soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_payload_we;
wire [26:0] soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_payload_addr;
reg soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_valid = 1'd0;
wire soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_ready;
reg soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_first = 1'd0;
reg soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_last = 1'd0;
reg [31:0] soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_payload_data = 32'd0;
reg soc_videooverlaysoc_out_dram_port_litedramnativeport1_flush = 1'd0;
reg soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_valid = 1'd0;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_ready;
reg soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_first = 1'd0;
reg soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_last = 1'd0;
reg [7:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_payload_sel = 8'd0;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_source_valid;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_source_ready;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_source_first;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_source_last;
wire [7:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_source_payload_sel;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_we;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_writable;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_re;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_readable;
wire [9:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_din;
wire [9:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_dout;
reg [2:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_level = 3'd0;
reg soc_videooverlaysoc_out_dram_port_cmd_buffer_replace = 1'd0;
reg [1:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_produce = 2'd0;
reg [1:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_consume = 2'd0;
reg [1:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_adr = 2'd0;
wire [9:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_dat_r;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_we;
wire [9:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_dat_w;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_do_read;
wire [1:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_rdport_adr;
wire [9:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_rdport_dat_r;
wire [7:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_in_payload_sel;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_in_first;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_in_last;
wire [7:0] soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_out_payload_sel;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_out_first;
wire soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_out_last;
reg [2:0] soc_videooverlaysoc_out_dram_port_counter = 3'd0;
reg soc_videooverlaysoc_out_dram_port_counter_ce = 1'd0;
wire soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_valid;
wire soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_ready;
wire soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_first;
wire soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_last;
wire [255:0] soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_payload_data;
wire soc_videooverlaysoc_out_dram_port_rdata_buffer_source_valid;
wire soc_videooverlaysoc_out_dram_port_rdata_buffer_source_ready;
wire soc_videooverlaysoc_out_dram_port_rdata_buffer_source_first;
wire soc_videooverlaysoc_out_dram_port_rdata_buffer_source_last;
reg [255:0] soc_videooverlaysoc_out_dram_port_rdata_buffer_source_payload_data = 256'd0;
wire soc_videooverlaysoc_out_dram_port_rdata_buffer_pipe_ce;
wire soc_videooverlaysoc_out_dram_port_rdata_buffer_busy;
reg soc_videooverlaysoc_out_dram_port_rdata_buffer_valid_n = 1'd0;
reg soc_videooverlaysoc_out_dram_port_rdata_buffer_first_n = 1'd0;
reg soc_videooverlaysoc_out_dram_port_rdata_buffer_last_n = 1'd0;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_sink_valid;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_sink_ready;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_sink_first;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_sink_last;
wire [255:0] soc_videooverlaysoc_out_dram_port_rdata_converter_sink_payload_data;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_source_valid;
reg soc_videooverlaysoc_out_dram_port_rdata_converter_source_ready = 1'd0;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_source_first;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_source_last;
wire [31:0] soc_videooverlaysoc_out_dram_port_rdata_converter_source_payload_data;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_valid;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_ready;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_first;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_last;
reg [255:0] soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data = 256'd0;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_valid;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_ready;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_first;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_last;
reg [31:0] soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data = 32'd0;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_valid_token_count;
reg [2:0] soc_videooverlaysoc_out_dram_port_rdata_converter_converter_mux = 3'd0;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_first;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_converter_last;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_valid;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_ready;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_first;
wire soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_last;
wire [31:0] soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_payload_data;
reg [7:0] soc_videooverlaysoc_out_dram_port_rdata_chunk = 8'd1;
wire soc_videooverlaysoc_out_dram_port_rdata_chunk_valid;
wire soc_videooverlaysoc_hdmi_core_out0_source_source_valid;
wire soc_videooverlaysoc_hdmi_core_out0_source_source_ready;
wire [23:0] soc_videooverlaysoc_hdmi_core_out0_source_source_payload_data;
wire soc_videooverlaysoc_hdmi_core_out0_source_source_param_hsync;
wire soc_videooverlaysoc_hdmi_core_out0_source_source_param_vsync;
wire soc_videooverlaysoc_hdmi_core_out0_source_source_param_de;
reg soc_videooverlaysoc_hdmi_core_out0_underflow_enable_storage_full = 1'd0;
wire soc_videooverlaysoc_hdmi_core_out0_underflow_enable_storage;
reg soc_videooverlaysoc_hdmi_core_out0_underflow_enable_re = 1'd0;
wire soc_videooverlaysoc_hdmi_core_out0_underflow_update_underflow_update_re;
wire soc_videooverlaysoc_hdmi_core_out0_underflow_update_underflow_update_r;
reg soc_videooverlaysoc_hdmi_core_out0_underflow_update_underflow_update_w = 1'd0;
reg [31:0] soc_videooverlaysoc_hdmi_core_out0_underflow_counter_status = 32'd0;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_valid;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_ready;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_first;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_last;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hscan;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vscan;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_base;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_length;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_valid;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_ready;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_first = 1'd0;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_last = 1'd0;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hscan;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vscan;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_base;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_length;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_valid;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_ready;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_first;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_last;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hscan;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vscan;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_base;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_length;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_we;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_writable;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_re;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_readable;
wire [161:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_din;
wire [161:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_dout;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [1:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q = 2'd0;
wire [1:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_next;
reg [1:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_binary = 2'd0;
reg [1:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_next_binary = 2'd0;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [1:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q = 2'd0;
wire [1:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next;
reg [1:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_binary = 2'd0;
reg [1:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next_binary = 2'd0;
wire [1:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_produce_rdomain;
wire [1:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_consume_wdomain;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_adr;
wire [161:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_dat_r;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_we;
wire [161:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_dat_w;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_rdport_adr;
wire [161:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_rdport_dat_r;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hscan;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vscan;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_base;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_length;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_first;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_last;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hscan;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vscan;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_base;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_length;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_first;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_last;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_enable_storage_full = 1'd0;
wire soc_videooverlaysoc_hdmi_core_out0_initiator_enable_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_enable_re = 1'd0;
reg [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_re = 1'd0;
reg [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_re = 1'd0;
reg [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_re = 1'd0;
reg [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_re = 1'd0;
reg [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_re = 1'd0;
reg [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_re = 1'd0;
reg [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_re = 1'd0;
reg [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_re = 1'd0;
reg [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage_full = 32'd0;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_re = 1'd0;
reg [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage_full = 32'd0;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage;
reg soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_re = 1'd0;
wire soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_valid;
reg soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_ready = 1'd0;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_hres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_hsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_hsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_hscan;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_vres;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_vsync_start;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_vsync_end;
wire [11:0] soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_vscan;
wire soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_valid;
reg soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_ready = 1'd0;
wire soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_first;
wire soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_last;
wire soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_hsync;
wire soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_vsync;
wire soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_de;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_valid;
reg soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_ready = 1'd0;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_payload_base;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_payload_length;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_source_valid;
reg soc_videooverlaysoc_hdmi_core_out0_dmareader_source_ready = 1'd0;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_source_first;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_source_last;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_source_payload_data;
reg soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_sink_valid = 1'd0;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_sink_ready;
wire [26:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_sink_payload_address;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_valid;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_ready;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_first;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_last;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_payload_data;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_request_enable;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_request_issued;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_data_dequeued;
reg [10:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_rsv_level = 11'd0;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_valid;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_ready;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_first;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_last;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_payload_data;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_valid;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_ready;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_first;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_last;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_payload_data;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_re;
reg soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_readable = 1'd0;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_we;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_writable;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_re;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_readable;
wire [33:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_din;
wire [33:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_dout;
reg [10:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level0 = 11'd0;
reg soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_replace = 1'd0;
reg [9:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_produce = 10'd0;
reg [9:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_consume = 10'd0;
reg [9:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_adr = 10'd0;
wire [33:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_dat_r;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_we;
wire [33:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_dat_w;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_do_read;
wire [9:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_rdport_adr;
wire [33:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_rdport_dat_r;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_rdport_re;
wire [10:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level1;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_in_payload_data;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_in_first;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_in_last;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_out_payload_data;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_out_first;
wire soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_out_last;
wire [26:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_base;
wire [26:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_length;
reg [26:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_offset = 27'd0;
reg [31:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full = 32'd0;
wire [31:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_storage;
reg soc_videooverlaysoc_hdmi_core_out0_dmareader_re = 1'd0;
reg soc_videooverlaysoc_hdmi_core_out0_dmareader_v = 1'd0;
reg soc_videooverlaysoc_hdmi_core_out0_dmareader_v_r = 1'd0;
reg soc_videooverlaysoc_hdmi_core_out0_dmareader_sof = 1'd0;
wire soc_videooverlaysoc_hdmi_core_out0_underflow_enable;
wire soc_videooverlaysoc_hdmi_core_out0_underflow_update;
reg [31:0] soc_videooverlaysoc_hdmi_core_out0_underflow_counter = 32'd0;
wire soc_videooverlaysoc_hdmi_core_out0_i;
wire soc_videooverlaysoc_hdmi_core_out0_o;
reg soc_videooverlaysoc_hdmi_core_out0_toggle_i = 1'd0;
wire soc_videooverlaysoc_hdmi_core_out0_toggle_o;
reg soc_videooverlaysoc_hdmi_core_out0_toggle_o_r = 1'd0;
reg soc_videooverlaysoc_core_source_valid_d = 1'd0;
reg [31:0] soc_videooverlaysoc_core_source_data_d = 32'd0;
wire soc_videooverlaysoc_timing_rgb_delay_sink_valid;
wire soc_videooverlaysoc_timing_rgb_delay_sink_ready;
wire soc_videooverlaysoc_timing_rgb_delay_sink_first;
wire soc_videooverlaysoc_timing_rgb_delay_sink_last;
wire [7:0] soc_videooverlaysoc_timing_rgb_delay_sink_payload_r;
wire [7:0] soc_videooverlaysoc_timing_rgb_delay_sink_payload_g;
wire [7:0] soc_videooverlaysoc_timing_rgb_delay_sink_payload_b;
reg soc_videooverlaysoc_timing_rgb_delay_source_valid = 1'd0;
reg soc_videooverlaysoc_timing_rgb_delay_source_ready = 1'd0;
reg soc_videooverlaysoc_timing_rgb_delay_source_first = 1'd0;
reg soc_videooverlaysoc_timing_rgb_delay_source_last = 1'd0;
wire [7:0] soc_videooverlaysoc_timing_rgb_delay_source_payload_r;
wire [7:0] soc_videooverlaysoc_timing_rgb_delay_source_payload_g;
wire [7:0] soc_videooverlaysoc_timing_rgb_delay_source_payload_b;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s0 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s1 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s2 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s3 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s4 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s5 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s6 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s7 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s8 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s9 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s10 = 8'd0;
reg [7:0] soc_videooverlaysoc_timing_rgb_delay_next_s11 = 8'd0;
wire soc_videooverlaysoc_hdmi_out0_rgb_valid;
reg soc_videooverlaysoc_hdmi_out0_rgb_ready = 1'd0;
reg soc_videooverlaysoc_hdmi_out0_rgb_first = 1'd0;
reg soc_videooverlaysoc_hdmi_out0_rgb_last = 1'd0;
wire [7:0] soc_videooverlaysoc_hdmi_out0_rgb_payload_r;
wire [7:0] soc_videooverlaysoc_hdmi_out0_rgb_payload_g;
wire [7:0] soc_videooverlaysoc_hdmi_out0_rgb_payload_b;
wire soc_videooverlaysoc_hdmi_out0_rgb_d_valid;
wire soc_videooverlaysoc_hdmi_out0_rgb_d_ready;
wire soc_videooverlaysoc_hdmi_out0_rgb_d_first;
wire soc_videooverlaysoc_hdmi_out0_rgb_d_last;
wire [7:0] soc_videooverlaysoc_hdmi_out0_rgb_d_payload_r;
wire [7:0] soc_videooverlaysoc_hdmi_out0_rgb_d_payload_g;
wire [7:0] soc_videooverlaysoc_hdmi_out0_rgb_d_payload_b;
reg [7:0] soc_videooverlaysoc_i2c_snoop_storage_full = 8'd0;
wire [7:0] soc_videooverlaysoc_i2c_snoop_storage;
reg soc_videooverlaysoc_i2c_snoop_re = 1'd0;
wire [7:0] soc_videooverlaysoc_i2c_snoop_status;
wire [7:0] soc_videooverlaysoc_i2c_snoop_reg_dout;
wire [63:0] soc_videooverlaysoc_i2c_snoop_An;
wire soc_videooverlaysoc_i2c_snoop_Aksv14_write;
wire soc_videooverlaysoc_hdcp_line_end;
reg soc_videooverlaysoc_hdcp_hpd = 1'd0;
reg soc_videooverlaysoc_hdcp_hdcp_ena = 1'd0;
reg soc_videooverlaysoc_hdcp_Aksv14_write = 1'd0;
reg [3:0] soc_videooverlaysoc_hdcp_ctl_code = 4'd0;
reg [63:0] soc_videooverlaysoc_hdcp_An = 64'd0;
reg [55:0] soc_videooverlaysoc_hdcp_Km_storage_full = 56'd0;
wire [55:0] soc_videooverlaysoc_hdcp_Km_storage;
reg soc_videooverlaysoc_hdcp_Km_re = 1'd0;
reg soc_videooverlaysoc_hdcp_Km_valid_storage_full = 1'd0;
wire soc_videooverlaysoc_hdcp_Km_valid_storage;
reg soc_videooverlaysoc_hdcp_Km_valid_re = 1'd0;
reg soc_videooverlaysoc_hdcp_hpd_ena_storage_full = 1'd0;
wire soc_videooverlaysoc_hdcp_hpd_ena_storage;
reg soc_videooverlaysoc_hdcp_hpd_ena_re = 1'd0;
wire [23:0] soc_videooverlaysoc_hdcp_cipher_stream;
wire soc_videooverlaysoc_hdcp_stream_ready;
wire soc_videooverlaysoc_Aksv14;
reg soc_videooverlaysoc_Aksv14_r = 1'd0;
reg [7:0] soc_videooverlaysoc_encoder0_d0 = 8'd0;
wire [1:0] soc_videooverlaysoc_encoder0_c;
wire soc_videooverlaysoc_encoder0_de;
reg [9:0] soc_videooverlaysoc_encoder0_out = 10'd0;
reg [7:0] soc_videooverlaysoc_encoder0_d1 = 8'd0;
reg [3:0] soc_videooverlaysoc_encoder0_n1d = 4'd0;
reg [8:0] soc_videooverlaysoc_encoder0_q_m = 9'd0;
wire soc_videooverlaysoc_encoder0_q_m8_n;
reg [8:0] soc_videooverlaysoc_encoder0_q_m_r = 9'd0;
reg [3:0] soc_videooverlaysoc_encoder0_n0q_m = 4'd0;
reg [3:0] soc_videooverlaysoc_encoder0_n1q_m = 4'd0;
reg signed [5:0] soc_videooverlaysoc_encoder0_cnt = 6'sd64;
reg [1:0] soc_videooverlaysoc_encoder0_new_c0 = 2'd0;
reg soc_videooverlaysoc_encoder0_new_de0 = 1'd0;
reg [1:0] soc_videooverlaysoc_encoder0_new_c1 = 2'd0;
reg soc_videooverlaysoc_encoder0_new_de1 = 1'd0;
reg [1:0] soc_videooverlaysoc_encoder0_new_c2 = 2'd0;
reg soc_videooverlaysoc_encoder0_new_de2 = 1'd0;
reg [7:0] soc_videooverlaysoc_encoder1_d0 = 8'd0;
wire [1:0] soc_videooverlaysoc_encoder1_c;
wire soc_videooverlaysoc_encoder1_de;
reg [9:0] soc_videooverlaysoc_encoder1_out = 10'd0;
reg [7:0] soc_videooverlaysoc_encoder1_d1 = 8'd0;
reg [3:0] soc_videooverlaysoc_encoder1_n1d = 4'd0;
reg [8:0] soc_videooverlaysoc_encoder1_q_m = 9'd0;
wire soc_videooverlaysoc_encoder1_q_m8_n;
reg [8:0] soc_videooverlaysoc_encoder1_q_m_r = 9'd0;
reg [3:0] soc_videooverlaysoc_encoder1_n0q_m = 4'd0;
reg [3:0] soc_videooverlaysoc_encoder1_n1q_m = 4'd0;
reg signed [5:0] soc_videooverlaysoc_encoder1_cnt = 6'sd64;
reg [1:0] soc_videooverlaysoc_encoder1_new_c0 = 2'd0;
reg soc_videooverlaysoc_encoder1_new_de0 = 1'd0;
reg [1:0] soc_videooverlaysoc_encoder1_new_c1 = 2'd0;
reg soc_videooverlaysoc_encoder1_new_de1 = 1'd0;
reg [1:0] soc_videooverlaysoc_encoder1_new_c2 = 2'd0;
reg soc_videooverlaysoc_encoder1_new_de2 = 1'd0;
reg [7:0] soc_videooverlaysoc_encoder2_d0 = 8'd0;
wire [1:0] soc_videooverlaysoc_encoder2_c;
wire soc_videooverlaysoc_encoder2_de;
reg [9:0] soc_videooverlaysoc_encoder2_out = 10'd0;
reg [7:0] soc_videooverlaysoc_encoder2_d1 = 8'd0;
reg [3:0] soc_videooverlaysoc_encoder2_n1d = 4'd0;
reg [8:0] soc_videooverlaysoc_encoder2_q_m = 9'd0;
wire soc_videooverlaysoc_encoder2_q_m8_n;
reg [8:0] soc_videooverlaysoc_encoder2_q_m_r = 9'd0;
reg [3:0] soc_videooverlaysoc_encoder2_n0q_m = 4'd0;
reg [3:0] soc_videooverlaysoc_encoder2_n1q_m = 4'd0;
reg signed [5:0] soc_videooverlaysoc_encoder2_cnt = 6'sd64;
reg [1:0] soc_videooverlaysoc_encoder2_new_c0 = 2'd0;
reg soc_videooverlaysoc_encoder2_new_de0 = 1'd0;
reg [1:0] soc_videooverlaysoc_encoder2_new_c1 = 2'd0;
reg soc_videooverlaysoc_encoder2_new_de1 = 1'd0;
reg [1:0] soc_videooverlaysoc_encoder2_new_c2 = 2'd0;
reg soc_videooverlaysoc_encoder2_new_de2 = 1'd0;
reg [9:0] soc_videooverlaysoc_c0_pix_o = 10'd0;
reg [9:0] soc_videooverlaysoc_c1_pix_o = 10'd0;
reg [9:0] soc_videooverlaysoc_c2_pix_o = 10'd0;
wire [9:0] soc_videooverlaysoc_c0;
wire [9:0] soc_videooverlaysoc_c1;
wire [9:0] soc_videooverlaysoc_c2;
reg [9:0] soc_videooverlaysoc_c0_next0 = 10'd0;
reg [9:0] soc_videooverlaysoc_c1_next0 = 10'd0;
reg [9:0] soc_videooverlaysoc_c2_next0 = 10'd0;
reg [9:0] soc_videooverlaysoc_c0_next1 = 10'd0;
reg [9:0] soc_videooverlaysoc_c1_next1 = 10'd0;
reg [9:0] soc_videooverlaysoc_c2_next1 = 10'd0;
reg [9:0] soc_videooverlaysoc_c0_next2 = 10'd0;
reg [9:0] soc_videooverlaysoc_c1_next2 = 10'd0;
reg [9:0] soc_videooverlaysoc_c2_next2 = 10'd0;
reg [9:0] soc_videooverlaysoc_c0_next3 = 10'd0;
reg [9:0] soc_videooverlaysoc_c1_next3 = 10'd0;
reg [9:0] soc_videooverlaysoc_c2_next3 = 10'd0;
reg [9:0] soc_videooverlaysoc_c0_next4 = 10'd0;
reg [9:0] soc_videooverlaysoc_c1_next4 = 10'd0;
reg [9:0] soc_videooverlaysoc_c2_next4 = 10'd0;
reg [9:0] soc_videooverlaysoc_c0_next5 = 10'd0;
reg [9:0] soc_videooverlaysoc_c1_next5 = 10'd0;
reg [9:0] soc_videooverlaysoc_c2_next5 = 10'd0;
wire soc_videooverlaysoc_rect_on0;
wire [7:0] soc_videooverlaysoc_rect_thresh;
reg [11:0] soc_videooverlaysoc_hrect_start_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_hrect_start_storage;
reg soc_videooverlaysoc_hrect_start_re = 1'd0;
reg [11:0] soc_videooverlaysoc_hrect_end_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_hrect_end_storage;
reg soc_videooverlaysoc_hrect_end_re = 1'd0;
reg [11:0] soc_videooverlaysoc_vrect_start_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_vrect_start_storage;
reg soc_videooverlaysoc_vrect_start_re = 1'd0;
reg [11:0] soc_videooverlaysoc_vrect_end_storage_full = 12'd0;
wire [11:0] soc_videooverlaysoc_vrect_end_storage;
reg soc_videooverlaysoc_vrect_end_re = 1'd0;
reg [7:0] soc_videooverlaysoc_rect_thresh_storage_full = 8'd0;
wire [7:0] soc_videooverlaysoc_rect_thresh_storage;
reg soc_videooverlaysoc_rect_thresh_re = 1'd0;
wire soc_videooverlaysoc_rect_on1;
reg [11:0] soc_videooverlaysoc_hcounter = 12'd0;
reg [11:0] soc_videooverlaysoc_vcounter = 12'd0;
reg soc_videooverlaysoc_in0_de = 1'd0;
reg soc_videooverlaysoc_in0_de_r = 1'd0;
reg soc_videooverlaysoc_in0_vsync = 1'd0;
reg soc_videooverlaysoc_in0_vsync_r = 1'd0;
reg soc_videooverlaysoc_in0_hsync = 1'd0;
reg soc_videooverlaysoc_in0_hsync_r = 1'd0;
reg soc_videooverlaysoc_phy_reset_storage = 1'd0;
wire eth_rx_clk;
wire eth_rx_rst;
wire eth_tx_clk;
wire eth_tx_rst;
wire soc_videooverlaysoc_phy_reset0;
wire soc_videooverlaysoc_phy_reset1;
reg [8:0] soc_videooverlaysoc_phy_counter = 9'd0;
wire soc_videooverlaysoc_phy_counter_done;
wire soc_videooverlaysoc_phy_counter_ce;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_ready;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_first;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_last;
wire [7:0] soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_payload_data;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_payload_last_be;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_payload_error;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_ready;
reg soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_first = 1'd0;
reg soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_last = 1'd0;
wire [7:0] soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_payload_data;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_ready;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_first;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_last;
wire [1:0] soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_payload_data;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_ready;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_first;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_last;
reg [7:0] soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_payload_data = 8'd0;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_ready;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_first;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_last;
reg [1:0] soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_payload_data = 2'd0;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_payload_valid_token_count;
reg [1:0] soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_mux = 2'd0;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_first;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_last;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_ready;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_first;
wire soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_last;
wire [1:0] soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_payload_data;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_ready;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_first;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_last;
wire [7:0] soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_payload_data;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_payload_last_be = 1'd0;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_payload_error = 1'd0;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_valid0;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_ready;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_first = 1'd0;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_last = 1'd0;
wire [1:0] soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_payload_data;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_ready;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_first;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_last;
reg [7:0] soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_payload_data = 8'd0;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_ready;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_first;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_last;
wire [1:0] soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_payload_data;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_ready;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_first = 1'd0;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_data = 8'd0;
reg [2:0] soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_valid_token_count = 3'd0;
reg [1:0] soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_demux = 2'd0;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_load_part;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_strobe_all = 1'd0;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_valid;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_ready;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_first;
wire soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_last;
wire [7:0] soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_payload_data;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_converter_reset = 1'd0;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_valid1 = 1'd0;
reg [1:0] soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_data = 2'd0;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_crs_dv = 1'd0;
reg soc_videooverlaysoc_phy_liteethphyrmiirx_crs_dv_d = 1'd0;
reg [1:0] soc_videooverlaysoc_phy_liteethphyrmiirx_rx_data = 2'd0;
reg [2:0] soc_videooverlaysoc_phy_storage = 3'd0;
wire soc_videooverlaysoc_phy_status;
wire soc_videooverlaysoc_phy_data_w;
wire soc_videooverlaysoc_phy_data_oe;
wire soc_videooverlaysoc_phy_data_r;
wire soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_valid;
reg soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_first;
wire soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_payload_data;
wire soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_payload_error;
reg soc_videooverlaysoc_core_mac_tx_gap_inserter_source_valid = 1'd0;
wire soc_videooverlaysoc_core_mac_tx_gap_inserter_source_ready;
reg soc_videooverlaysoc_core_mac_tx_gap_inserter_source_first = 1'd0;
reg soc_videooverlaysoc_core_mac_tx_gap_inserter_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_last_be = 1'd0;
reg soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_error = 1'd0;
reg [3:0] soc_videooverlaysoc_core_mac_tx_gap_inserter_counter = 4'd0;
reg soc_videooverlaysoc_core_mac_tx_gap_inserter_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_mac_tx_gap_inserter_counter_ce = 1'd0;
reg [31:0] soc_videooverlaysoc_core_mac_preamble_errors_status = 32'd0;
reg [31:0] soc_videooverlaysoc_core_mac_crc_errors_status = 32'd0;
wire soc_videooverlaysoc_core_mac_preamble_inserter_sink_valid;
reg soc_videooverlaysoc_core_mac_preamble_inserter_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_mac_preamble_inserter_sink_first;
wire soc_videooverlaysoc_core_mac_preamble_inserter_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_preamble_inserter_sink_payload_data;
wire soc_videooverlaysoc_core_mac_preamble_inserter_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_preamble_inserter_sink_payload_error;
reg soc_videooverlaysoc_core_mac_preamble_inserter_source_valid = 1'd0;
wire soc_videooverlaysoc_core_mac_preamble_inserter_source_ready;
reg soc_videooverlaysoc_core_mac_preamble_inserter_source_first = 1'd0;
reg soc_videooverlaysoc_core_mac_preamble_inserter_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data = 8'd0;
wire soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_last_be;
reg soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_error = 1'd0;
reg [63:0] soc_videooverlaysoc_core_mac_preamble_inserter_preamble = 64'd15372286728091293013;
reg [2:0] soc_videooverlaysoc_core_mac_preamble_inserter_cnt = 3'd0;
reg soc_videooverlaysoc_core_mac_preamble_inserter_clr_cnt = 1'd0;
reg soc_videooverlaysoc_core_mac_preamble_inserter_inc_cnt = 1'd0;
wire soc_videooverlaysoc_core_mac_preamble_checker_sink_valid;
reg soc_videooverlaysoc_core_mac_preamble_checker_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_mac_preamble_checker_sink_first;
wire soc_videooverlaysoc_core_mac_preamble_checker_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_preamble_checker_sink_payload_data;
wire soc_videooverlaysoc_core_mac_preamble_checker_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_preamble_checker_sink_payload_error;
reg soc_videooverlaysoc_core_mac_preamble_checker_source_valid = 1'd0;
wire soc_videooverlaysoc_core_mac_preamble_checker_source_ready;
reg soc_videooverlaysoc_core_mac_preamble_checker_source_first = 1'd0;
reg soc_videooverlaysoc_core_mac_preamble_checker_source_last = 1'd0;
wire [7:0] soc_videooverlaysoc_core_mac_preamble_checker_source_payload_data;
wire soc_videooverlaysoc_core_mac_preamble_checker_source_payload_last_be;
reg soc_videooverlaysoc_core_mac_preamble_checker_source_payload_error = 1'd0;
reg soc_videooverlaysoc_core_mac_preamble_checker_error = 1'd0;
wire soc_videooverlaysoc_core_mac_crc32_inserter_sink_valid;
reg soc_videooverlaysoc_core_mac_crc32_inserter_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_mac_crc32_inserter_sink_first;
wire soc_videooverlaysoc_core_mac_crc32_inserter_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_crc32_inserter_sink_payload_data;
wire soc_videooverlaysoc_core_mac_crc32_inserter_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_crc32_inserter_sink_payload_error;
reg soc_videooverlaysoc_core_mac_crc32_inserter_source_valid = 1'd0;
wire soc_videooverlaysoc_core_mac_crc32_inserter_source_ready;
reg soc_videooverlaysoc_core_mac_crc32_inserter_source_first = 1'd0;
reg soc_videooverlaysoc_core_mac_crc32_inserter_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_last_be = 1'd0;
reg soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_error = 1'd0;
reg [7:0] soc_videooverlaysoc_core_mac_crc32_inserter_data0 = 8'd0;
wire [31:0] soc_videooverlaysoc_core_mac_crc32_inserter_value;
wire soc_videooverlaysoc_core_mac_crc32_inserter_error;
wire [7:0] soc_videooverlaysoc_core_mac_crc32_inserter_data1;
wire [31:0] soc_videooverlaysoc_core_mac_crc32_inserter_last;
reg [31:0] soc_videooverlaysoc_core_mac_crc32_inserter_next = 32'd0;
reg [31:0] soc_videooverlaysoc_core_mac_crc32_inserter_reg = 32'd4294967295;
reg soc_videooverlaysoc_core_mac_crc32_inserter_ce = 1'd0;
reg soc_videooverlaysoc_core_mac_crc32_inserter_reset = 1'd0;
reg [1:0] soc_videooverlaysoc_core_mac_crc32_inserter_cnt = 2'd3;
wire soc_videooverlaysoc_core_mac_crc32_inserter_cnt_done;
reg soc_videooverlaysoc_core_mac_crc32_inserter_is_ongoing0 = 1'd0;
reg soc_videooverlaysoc_core_mac_crc32_inserter_is_ongoing1 = 1'd0;
wire soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_valid;
reg soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_first;
wire soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_data;
wire soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_error;
wire soc_videooverlaysoc_core_mac_crc32_checker_source_source_valid;
wire soc_videooverlaysoc_core_mac_crc32_checker_source_source_ready;
reg soc_videooverlaysoc_core_mac_crc32_checker_source_source_first = 1'd0;
wire soc_videooverlaysoc_core_mac_crc32_checker_source_source_last;
wire [7:0] soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_data;
wire soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_last_be;
reg soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_error = 1'd0;
wire soc_videooverlaysoc_core_mac_crc32_checker_error;
wire [7:0] soc_videooverlaysoc_core_mac_crc32_checker_crc_data0;
wire [31:0] soc_videooverlaysoc_core_mac_crc32_checker_crc_value;
wire soc_videooverlaysoc_core_mac_crc32_checker_crc_error;
wire [7:0] soc_videooverlaysoc_core_mac_crc32_checker_crc_data1;
wire [31:0] soc_videooverlaysoc_core_mac_crc32_checker_crc_last;
reg [31:0] soc_videooverlaysoc_core_mac_crc32_checker_crc_next = 32'd0;
reg [31:0] soc_videooverlaysoc_core_mac_crc32_checker_crc_reg = 32'd4294967295;
reg soc_videooverlaysoc_core_mac_crc32_checker_crc_ce = 1'd0;
reg soc_videooverlaysoc_core_mac_crc32_checker_crc_reset = 1'd0;
reg soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_valid = 1'd0;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_ready;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_first;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_payload_data;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_payload_error;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_valid;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_ready;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_first;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_last;
wire [7:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_payload_data;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_payload_last_be;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_payload_error;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_we;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_writable;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_re;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_readable;
wire [11:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_din;
wire [11:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_dout;
reg [2:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_level = 3'd0;
reg soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_replace = 1'd0;
reg [2:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_produce = 3'd0;
reg [2:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_consume = 3'd0;
reg [2:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_adr = 3'd0;
wire [11:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_dat_r;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_we;
wire [11:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_dat_w;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_do_read;
wire [2:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_rdport_adr;
wire [11:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_rdport_dat_r;
wire [7:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_payload_data;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_payload_last_be;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_payload_error;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_first;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_last;
wire [7:0] soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_payload_data;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_payload_last_be;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_payload_error;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_first;
wire soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_last;
reg soc_videooverlaysoc_core_mac_crc32_checker_fifo_reset = 1'd0;
wire soc_videooverlaysoc_core_mac_crc32_checker_fifo_in;
wire soc_videooverlaysoc_core_mac_crc32_checker_fifo_out;
wire soc_videooverlaysoc_core_mac_crc32_checker_fifo_full;
wire soc_videooverlaysoc_core_mac_ps_preamble_error_i;
wire soc_videooverlaysoc_core_mac_ps_preamble_error_o;
reg soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_i = 1'd0;
wire soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_o;
reg soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_core_mac_ps_crc_error_i;
wire soc_videooverlaysoc_core_mac_ps_crc_error_o;
reg soc_videooverlaysoc_core_mac_ps_crc_error_toggle_i = 1'd0;
wire soc_videooverlaysoc_core_mac_ps_crc_error_toggle_o;
reg soc_videooverlaysoc_core_mac_ps_crc_error_toggle_o_r = 1'd0;
wire soc_videooverlaysoc_core_mac_padding_inserter_sink_valid;
reg soc_videooverlaysoc_core_mac_padding_inserter_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_mac_padding_inserter_sink_first;
wire soc_videooverlaysoc_core_mac_padding_inserter_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_padding_inserter_sink_payload_data;
wire soc_videooverlaysoc_core_mac_padding_inserter_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_padding_inserter_sink_payload_error;
reg soc_videooverlaysoc_core_mac_padding_inserter_source_valid = 1'd0;
wire soc_videooverlaysoc_core_mac_padding_inserter_source_ready;
reg soc_videooverlaysoc_core_mac_padding_inserter_source_first = 1'd0;
reg soc_videooverlaysoc_core_mac_padding_inserter_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_mac_padding_inserter_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_mac_padding_inserter_source_payload_last_be = 1'd0;
reg soc_videooverlaysoc_core_mac_padding_inserter_source_payload_error = 1'd0;
reg [15:0] soc_videooverlaysoc_core_mac_padding_inserter_counter = 16'd1;
wire soc_videooverlaysoc_core_mac_padding_inserter_counter_done;
reg soc_videooverlaysoc_core_mac_padding_inserter_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_mac_padding_inserter_counter_ce = 1'd0;
wire soc_videooverlaysoc_core_mac_padding_checker_sink_valid;
wire soc_videooverlaysoc_core_mac_padding_checker_sink_ready;
wire soc_videooverlaysoc_core_mac_padding_checker_sink_first;
wire soc_videooverlaysoc_core_mac_padding_checker_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_padding_checker_sink_payload_data;
wire soc_videooverlaysoc_core_mac_padding_checker_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_padding_checker_sink_payload_error;
wire soc_videooverlaysoc_core_mac_padding_checker_source_valid;
wire soc_videooverlaysoc_core_mac_padding_checker_source_ready;
wire soc_videooverlaysoc_core_mac_padding_checker_source_first;
wire soc_videooverlaysoc_core_mac_padding_checker_source_last;
wire [7:0] soc_videooverlaysoc_core_mac_padding_checker_source_payload_data;
wire soc_videooverlaysoc_core_mac_padding_checker_source_payload_last_be;
wire soc_videooverlaysoc_core_mac_padding_checker_source_payload_error;
wire soc_videooverlaysoc_core_mac_tx_cdc_sink_valid;
wire soc_videooverlaysoc_core_mac_tx_cdc_sink_ready;
wire soc_videooverlaysoc_core_mac_tx_cdc_sink_first;
wire soc_videooverlaysoc_core_mac_tx_cdc_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_tx_cdc_sink_payload_data;
wire soc_videooverlaysoc_core_mac_tx_cdc_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_tx_cdc_sink_payload_error;
wire soc_videooverlaysoc_core_mac_tx_cdc_source_valid;
wire soc_videooverlaysoc_core_mac_tx_cdc_source_ready;
wire soc_videooverlaysoc_core_mac_tx_cdc_source_first;
wire soc_videooverlaysoc_core_mac_tx_cdc_source_last;
wire [7:0] soc_videooverlaysoc_core_mac_tx_cdc_source_payload_data;
wire soc_videooverlaysoc_core_mac_tx_cdc_source_payload_last_be;
wire soc_videooverlaysoc_core_mac_tx_cdc_source_payload_error;
wire soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_we;
wire soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_writable;
wire soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_re;
wire soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_readable;
wire [11:0] soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_din;
wire [11:0] soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_dout;
wire soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q = 7'd0;
wire [6:0] soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_next;
reg [6:0] soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_next_binary = 7'd0;
wire soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q = 7'd0;
wire [6:0] soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next;
reg [6:0] soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next_binary = 7'd0;
wire [6:0] soc_videooverlaysoc_core_mac_tx_cdc_produce_rdomain;
wire [6:0] soc_videooverlaysoc_core_mac_tx_cdc_consume_wdomain;
wire [5:0] soc_videooverlaysoc_core_mac_tx_cdc_wrport_adr;
wire [11:0] soc_videooverlaysoc_core_mac_tx_cdc_wrport_dat_r;
wire soc_videooverlaysoc_core_mac_tx_cdc_wrport_we;
wire [11:0] soc_videooverlaysoc_core_mac_tx_cdc_wrport_dat_w;
wire [5:0] soc_videooverlaysoc_core_mac_tx_cdc_rdport_adr;
wire [11:0] soc_videooverlaysoc_core_mac_tx_cdc_rdport_dat_r;
wire [7:0] soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_payload_data;
wire soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_payload_last_be;
wire soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_payload_error;
wire soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_first;
wire soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_last;
wire [7:0] soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_payload_data;
wire soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_payload_last_be;
wire soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_payload_error;
wire soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_first;
wire soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_last;
wire soc_videooverlaysoc_core_mac_rx_cdc_sink_valid;
wire soc_videooverlaysoc_core_mac_rx_cdc_sink_ready;
wire soc_videooverlaysoc_core_mac_rx_cdc_sink_first;
wire soc_videooverlaysoc_core_mac_rx_cdc_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_rx_cdc_sink_payload_data;
wire soc_videooverlaysoc_core_mac_rx_cdc_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_rx_cdc_sink_payload_error;
wire soc_videooverlaysoc_core_mac_rx_cdc_source_valid;
wire soc_videooverlaysoc_core_mac_rx_cdc_source_ready;
wire soc_videooverlaysoc_core_mac_rx_cdc_source_first;
wire soc_videooverlaysoc_core_mac_rx_cdc_source_last;
wire [7:0] soc_videooverlaysoc_core_mac_rx_cdc_source_payload_data;
wire soc_videooverlaysoc_core_mac_rx_cdc_source_payload_last_be;
wire soc_videooverlaysoc_core_mac_rx_cdc_source_payload_error;
wire soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_we;
wire soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_writable;
wire soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_re;
wire soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_readable;
wire [11:0] soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_din;
wire [11:0] soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_dout;
wire soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q = 7'd0;
wire [6:0] soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_next;
reg [6:0] soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_next_binary = 7'd0;
wire soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q = 7'd0;
wire [6:0] soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next;
reg [6:0] soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next_binary = 7'd0;
wire [6:0] soc_videooverlaysoc_core_mac_rx_cdc_produce_rdomain;
wire [6:0] soc_videooverlaysoc_core_mac_rx_cdc_consume_wdomain;
wire [5:0] soc_videooverlaysoc_core_mac_rx_cdc_wrport_adr;
wire [11:0] soc_videooverlaysoc_core_mac_rx_cdc_wrport_dat_r;
wire soc_videooverlaysoc_core_mac_rx_cdc_wrport_we;
wire [11:0] soc_videooverlaysoc_core_mac_rx_cdc_wrport_dat_w;
wire [5:0] soc_videooverlaysoc_core_mac_rx_cdc_rdport_adr;
wire [11:0] soc_videooverlaysoc_core_mac_rx_cdc_rdport_dat_r;
wire [7:0] soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_payload_data;
wire soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_payload_last_be;
wire soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_payload_error;
wire soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_first;
wire soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_last;
wire [7:0] soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_payload_data;
wire soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_payload_last_be;
wire soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_payload_error;
wire soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_first;
wire soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_last;
reg soc_videooverlaysoc_core_mac_crossbar_source_valid = 1'd0;
wire soc_videooverlaysoc_core_mac_crossbar_source_ready;
reg soc_videooverlaysoc_core_mac_crossbar_source_first = 1'd0;
reg soc_videooverlaysoc_core_mac_crossbar_source_last = 1'd0;
reg [15:0] soc_videooverlaysoc_core_mac_crossbar_source_payload_ethernet_type = 16'd0;
reg [47:0] soc_videooverlaysoc_core_mac_crossbar_source_payload_sender_mac = 48'd0;
reg [47:0] soc_videooverlaysoc_core_mac_crossbar_source_payload_target_mac = 48'd0;
reg [7:0] soc_videooverlaysoc_core_mac_crossbar_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_mac_crossbar_source_payload_last_be = 1'd0;
reg soc_videooverlaysoc_core_mac_crossbar_source_payload_error = 1'd0;
wire soc_videooverlaysoc_core_mac_crossbar_sink_valid;
reg soc_videooverlaysoc_core_mac_crossbar_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_mac_crossbar_sink_first;
wire soc_videooverlaysoc_core_mac_crossbar_sink_last;
wire [15:0] soc_videooverlaysoc_core_mac_crossbar_sink_payload_ethernet_type;
wire [47:0] soc_videooverlaysoc_core_mac_crossbar_sink_payload_sender_mac;
wire [47:0] soc_videooverlaysoc_core_mac_crossbar_sink_payload_target_mac;
wire [7:0] soc_videooverlaysoc_core_mac_crossbar_sink_payload_data;
wire soc_videooverlaysoc_core_mac_crossbar_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_crossbar_sink_payload_error;
wire soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_valid;
reg soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_first;
wire soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_last;
wire [15:0] soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_ethernet_type;
wire [47:0] soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_sender_mac;
wire [47:0] soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_target_mac;
wire [7:0] soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_data;
wire soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_error;
reg soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_valid = 1'd0;
wire soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_ready;
reg soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_first = 1'd0;
reg soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_last_be = 1'd0;
wire soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_error;
reg [111:0] soc_videooverlaysoc_core_mac_liteethmacpacketizer_header = 112'd0;
reg [111:0] soc_videooverlaysoc_core_mac_liteethmacpacketizer_header_reg = 112'd0;
reg soc_videooverlaysoc_core_mac_liteethmacpacketizer_load = 1'd0;
reg soc_videooverlaysoc_core_mac_liteethmacpacketizer_shift = 1'd0;
reg [3:0] soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter = 4'd0;
reg soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter_ce = 1'd0;
reg [7:0] soc_videooverlaysoc_core_mac_liteethmacpacketizer = 8'd0;
wire soc_videooverlaysoc_core_mac_depacketizer_sink_valid;
reg soc_videooverlaysoc_core_mac_depacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_mac_depacketizer_sink_first;
wire soc_videooverlaysoc_core_mac_depacketizer_sink_last;
wire [7:0] soc_videooverlaysoc_core_mac_depacketizer_sink_payload_data;
wire soc_videooverlaysoc_core_mac_depacketizer_sink_payload_last_be;
wire soc_videooverlaysoc_core_mac_depacketizer_sink_payload_error;
reg soc_videooverlaysoc_core_mac_depacketizer_source_valid = 1'd0;
wire soc_videooverlaysoc_core_mac_depacketizer_source_ready;
reg soc_videooverlaysoc_core_mac_depacketizer_source_first = 1'd0;
wire soc_videooverlaysoc_core_mac_depacketizer_source_last;
wire [15:0] soc_videooverlaysoc_core_mac_depacketizer_source_payload_ethernet_type;
wire [47:0] soc_videooverlaysoc_core_mac_depacketizer_source_payload_sender_mac;
wire [47:0] soc_videooverlaysoc_core_mac_depacketizer_source_payload_target_mac;
wire [7:0] soc_videooverlaysoc_core_mac_depacketizer_source_payload_data;
reg soc_videooverlaysoc_core_mac_depacketizer_source_payload_last_be = 1'd0;
wire soc_videooverlaysoc_core_mac_depacketizer_source_payload_error;
wire [111:0] soc_videooverlaysoc_core_mac_depacketizer_header;
reg [111:0] soc_videooverlaysoc_core_mac_depacketizer_header_reg = 112'd0;
reg soc_videooverlaysoc_core_mac_depacketizer_shift = 1'd0;
reg [3:0] soc_videooverlaysoc_core_mac_depacketizer_counter = 4'd0;
reg soc_videooverlaysoc_core_mac_depacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_mac_depacketizer_counter_ce = 1'd0;
reg soc_videooverlaysoc_core_mac_depacketizer_no_payload = 1'd0;
wire soc_videooverlaysoc_core_mac_depacketizer_is_el;
wire soc_videooverlaysoc_core_arp_tx_sink_valid;
reg soc_videooverlaysoc_core_arp_tx_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_arp_tx_sink_first;
wire soc_videooverlaysoc_core_arp_tx_sink_last;
wire soc_videooverlaysoc_core_arp_tx_sink_payload_reply;
wire soc_videooverlaysoc_core_arp_tx_sink_payload_request;
wire [31:0] soc_videooverlaysoc_core_arp_tx_sink_payload_ip_address;
wire [47:0] soc_videooverlaysoc_core_arp_tx_sink_payload_mac_address;
reg soc_videooverlaysoc_core_arp_tx_source_valid = 1'd0;
wire soc_videooverlaysoc_core_arp_tx_source_ready;
reg soc_videooverlaysoc_core_arp_tx_source_first = 1'd0;
reg soc_videooverlaysoc_core_arp_tx_source_last = 1'd0;
reg [15:0] soc_videooverlaysoc_core_arp_tx_source_payload_ethernet_type = 16'd0;
reg [47:0] soc_videooverlaysoc_core_arp_tx_source_payload_sender_mac = 48'd0;
reg [47:0] soc_videooverlaysoc_core_arp_tx_source_payload_target_mac = 48'd0;
reg [7:0] soc_videooverlaysoc_core_arp_tx_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_arp_tx_source_payload_last_be = 1'd0;
reg soc_videooverlaysoc_core_arp_tx_source_payload_error = 1'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_valid = 1'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_last;
reg [7:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_payload_data = 8'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_payload_error = 1'd0;
wire [7:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_hwsize;
wire [15:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_hwtype;
reg [15:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_opcode = 16'd0;
wire [15:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_proto;
wire [7:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_protosize;
wire [31:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_ip;
wire [47:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_mac;
reg [31:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_ip = 32'd0;
reg [47:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac = 48'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_valid = 1'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_ready = 1'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_first = 1'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_last = 1'd0;
reg [15:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_ethernet_type = 16'd0;
reg [47:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_sender_mac = 48'd0;
reg [47:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_target_mac = 48'd0;
reg [7:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_last_be = 1'd0;
wire soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_error;
reg [223:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header = 224'd0;
reg [223:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header_reg = 224'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_load = 1'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_shift = 1'd0;
reg [4:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter = 5'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter_ce = 1'd0;
reg [7:0] soc_videooverlaysoc_core_arp_tx_liteetharppacketizer = 8'd0;
reg [5:0] soc_videooverlaysoc_core_arp_tx_counter = 6'd0;
reg soc_videooverlaysoc_core_arp_tx_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_arp_tx_counter_ce = 1'd0;
wire soc_videooverlaysoc_core_arp_sink_sink_valid;
wire soc_videooverlaysoc_core_arp_sink_sink_ready;
wire soc_videooverlaysoc_core_arp_sink_sink_first;
wire soc_videooverlaysoc_core_arp_sink_sink_last;
wire [15:0] soc_videooverlaysoc_core_arp_sink_sink_payload_ethernet_type;
wire [47:0] soc_videooverlaysoc_core_arp_sink_sink_payload_sender_mac;
wire [47:0] soc_videooverlaysoc_core_arp_sink_sink_payload_target_mac;
wire [7:0] soc_videooverlaysoc_core_arp_sink_sink_payload_data;
wire soc_videooverlaysoc_core_arp_sink_sink_payload_last_be;
wire soc_videooverlaysoc_core_arp_sink_sink_payload_error;
reg soc_videooverlaysoc_core_arp_source_source_valid = 1'd0;
wire soc_videooverlaysoc_core_arp_source_source_ready;
reg soc_videooverlaysoc_core_arp_source_source_first = 1'd0;
reg soc_videooverlaysoc_core_arp_source_source_last = 1'd0;
reg soc_videooverlaysoc_core_arp_source_source_payload_reply = 1'd0;
reg soc_videooverlaysoc_core_arp_source_source_payload_request = 1'd0;
wire [31:0] soc_videooverlaysoc_core_arp_source_source_payload_ip_address;
wire [47:0] soc_videooverlaysoc_core_arp_source_source_payload_mac_address;
wire soc_videooverlaysoc_core_arp_depacketizer_sink_valid;
reg soc_videooverlaysoc_core_arp_depacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_arp_depacketizer_sink_first;
wire soc_videooverlaysoc_core_arp_depacketizer_sink_last;
wire [15:0] soc_videooverlaysoc_core_arp_depacketizer_sink_payload_ethernet_type;
wire [47:0] soc_videooverlaysoc_core_arp_depacketizer_sink_payload_sender_mac;
wire [47:0] soc_videooverlaysoc_core_arp_depacketizer_sink_payload_target_mac;
wire [7:0] soc_videooverlaysoc_core_arp_depacketizer_sink_payload_data;
wire soc_videooverlaysoc_core_arp_depacketizer_sink_payload_last_be;
wire soc_videooverlaysoc_core_arp_depacketizer_sink_payload_error;
reg soc_videooverlaysoc_core_arp_depacketizer_source_valid = 1'd0;
reg soc_videooverlaysoc_core_arp_depacketizer_source_ready = 1'd0;
wire soc_videooverlaysoc_core_arp_depacketizer_source_last;
wire [7:0] soc_videooverlaysoc_core_arp_depacketizer_source_payload_data;
wire soc_videooverlaysoc_core_arp_depacketizer_source_payload_error;
wire [7:0] soc_videooverlaysoc_core_arp_depacketizer_source_param_hwsize;
wire [15:0] soc_videooverlaysoc_core_arp_depacketizer_source_param_hwtype;
wire [15:0] soc_videooverlaysoc_core_arp_depacketizer_source_param_opcode;
wire [15:0] soc_videooverlaysoc_core_arp_depacketizer_source_param_proto;
wire [7:0] soc_videooverlaysoc_core_arp_depacketizer_source_param_protosize;
wire [31:0] soc_videooverlaysoc_core_arp_depacketizer_source_param_sender_ip;
wire [47:0] soc_videooverlaysoc_core_arp_depacketizer_source_param_sender_mac;
wire [31:0] soc_videooverlaysoc_core_arp_depacketizer_source_param_target_ip;
wire [47:0] soc_videooverlaysoc_core_arp_depacketizer_source_param_target_mac;
wire [223:0] soc_videooverlaysoc_core_arp_depacketizer_header;
reg [223:0] soc_videooverlaysoc_core_arp_depacketizer_header_reg = 224'd0;
reg soc_videooverlaysoc_core_arp_depacketizer_shift = 1'd0;
reg [4:0] soc_videooverlaysoc_core_arp_depacketizer_counter = 5'd0;
reg soc_videooverlaysoc_core_arp_depacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_arp_depacketizer_counter_ce = 1'd0;
reg soc_videooverlaysoc_core_arp_depacketizer_no_payload = 1'd0;
wire soc_videooverlaysoc_core_arp_depacketizer_is_el;
reg soc_videooverlaysoc_core_arp_valid = 1'd0;
reg soc_videooverlaysoc_core_arp_reply = 1'd0;
reg soc_videooverlaysoc_core_arp_request = 1'd0;
wire soc_videooverlaysoc_core_arp_table_sink_valid;
reg soc_videooverlaysoc_core_arp_table_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_arp_table_sink_first;
wire soc_videooverlaysoc_core_arp_table_sink_last;
wire soc_videooverlaysoc_core_arp_table_sink_payload_reply;
wire soc_videooverlaysoc_core_arp_table_sink_payload_request;
wire [31:0] soc_videooverlaysoc_core_arp_table_sink_payload_ip_address;
wire [47:0] soc_videooverlaysoc_core_arp_table_sink_payload_mac_address;
reg soc_videooverlaysoc_core_arp_table_source_valid = 1'd0;
wire soc_videooverlaysoc_core_arp_table_source_ready;
reg soc_videooverlaysoc_core_arp_table_source_first = 1'd0;
reg soc_videooverlaysoc_core_arp_table_source_last = 1'd0;
reg soc_videooverlaysoc_core_arp_table_source_payload_reply = 1'd0;
reg soc_videooverlaysoc_core_arp_table_source_payload_request = 1'd0;
reg [31:0] soc_videooverlaysoc_core_arp_table_source_payload_ip_address = 32'd0;
reg [47:0] soc_videooverlaysoc_core_arp_table_source_payload_mac_address = 48'd0;
reg soc_videooverlaysoc_core_arp_table_request_valid = 1'd0;
reg soc_videooverlaysoc_core_arp_table_request_ready = 1'd0;
wire [31:0] soc_videooverlaysoc_core_arp_table_request_payload_ip_address;
reg soc_videooverlaysoc_core_arp_table_response_valid = 1'd0;
reg soc_videooverlaysoc_core_arp_table_response_ready = 1'd0;
reg soc_videooverlaysoc_core_arp_table_response_payload_failed = 1'd0;
wire [47:0] soc_videooverlaysoc_core_arp_table_response_payload_mac_address;
reg soc_videooverlaysoc_core_arp_table_request_pending = 1'd0;
reg soc_videooverlaysoc_core_arp_table_request_pending_clr = 1'd0;
reg soc_videooverlaysoc_core_arp_table_request_pending_set = 1'd0;
reg [31:0] soc_videooverlaysoc_core_arp_table_request_ip_address = 32'd0;
reg soc_videooverlaysoc_core_arp_table_request_ip_address_reset = 1'd0;
reg soc_videooverlaysoc_core_arp_table_request_ip_address_update = 1'd0;
wire soc_videooverlaysoc_core_arp_table_request_timer_wait;
wire soc_videooverlaysoc_core_arp_table_request_timer_done;
reg [22:0] soc_videooverlaysoc_core_arp_table_request_timer_count = 23'd5000000;
reg [2:0] soc_videooverlaysoc_core_arp_table_request_counter = 3'd0;
reg soc_videooverlaysoc_core_arp_table_request_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_arp_table_request_counter_ce = 1'd0;
reg soc_videooverlaysoc_core_arp_table_update = 1'd0;
reg soc_videooverlaysoc_core_arp_table_cached_valid = 1'd0;
reg [31:0] soc_videooverlaysoc_core_arp_table_cached_ip_address = 32'd0;
reg [47:0] soc_videooverlaysoc_core_arp_table_cached_mac_address = 48'd0;
wire soc_videooverlaysoc_core_arp_table_cached_timer_wait;
wire soc_videooverlaysoc_core_arp_table_cached_timer_done;
reg [28:0] soc_videooverlaysoc_core_arp_table_cached_timer_count = 29'd500000000;
wire soc_videooverlaysoc_core_arp_mac_port_sink_valid;
reg soc_videooverlaysoc_core_arp_mac_port_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_arp_mac_port_sink_first;
wire soc_videooverlaysoc_core_arp_mac_port_sink_last;
wire [15:0] soc_videooverlaysoc_core_arp_mac_port_sink_payload_ethernet_type;
wire [47:0] soc_videooverlaysoc_core_arp_mac_port_sink_payload_sender_mac;
wire [47:0] soc_videooverlaysoc_core_arp_mac_port_sink_payload_target_mac;
wire [7:0] soc_videooverlaysoc_core_arp_mac_port_sink_payload_data;
wire soc_videooverlaysoc_core_arp_mac_port_sink_payload_last_be;
wire soc_videooverlaysoc_core_arp_mac_port_sink_payload_error;
reg soc_videooverlaysoc_core_arp_mac_port_source_valid = 1'd0;
wire soc_videooverlaysoc_core_arp_mac_port_source_ready;
reg soc_videooverlaysoc_core_arp_mac_port_source_first = 1'd0;
reg soc_videooverlaysoc_core_arp_mac_port_source_last = 1'd0;
reg [15:0] soc_videooverlaysoc_core_arp_mac_port_source_payload_ethernet_type = 16'd0;
reg [47:0] soc_videooverlaysoc_core_arp_mac_port_source_payload_sender_mac = 48'd0;
reg [47:0] soc_videooverlaysoc_core_arp_mac_port_source_payload_target_mac = 48'd0;
reg [7:0] soc_videooverlaysoc_core_arp_mac_port_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_arp_mac_port_source_payload_last_be = 1'd0;
reg soc_videooverlaysoc_core_arp_mac_port_source_payload_error = 1'd0;
wire soc_videooverlaysoc_core_ip_tx_sink_valid;
wire soc_videooverlaysoc_core_ip_tx_sink_ready;
wire soc_videooverlaysoc_core_ip_tx_sink_first;
wire soc_videooverlaysoc_core_ip_tx_sink_last;
wire [7:0] soc_videooverlaysoc_core_ip_tx_sink_payload_data;
wire soc_videooverlaysoc_core_ip_tx_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_ip_tx_sink_param_length;
wire [7:0] soc_videooverlaysoc_core_ip_tx_sink_param_protocol;
wire [31:0] soc_videooverlaysoc_core_ip_tx_sink_param_ip_address;
reg soc_videooverlaysoc_core_ip_tx_source_valid = 1'd0;
wire soc_videooverlaysoc_core_ip_tx_source_ready;
reg soc_videooverlaysoc_core_ip_tx_source_first = 1'd0;
reg soc_videooverlaysoc_core_ip_tx_source_last = 1'd0;
reg [15:0] soc_videooverlaysoc_core_ip_tx_source_payload_ethernet_type = 16'd0;
reg [47:0] soc_videooverlaysoc_core_ip_tx_source_payload_sender_mac = 48'd0;
reg [47:0] soc_videooverlaysoc_core_ip_tx_source_payload_target_mac = 48'd0;
reg [7:0] soc_videooverlaysoc_core_ip_tx_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_ip_tx_source_payload_last_be = 1'd0;
reg soc_videooverlaysoc_core_ip_tx_source_payload_error = 1'd0;
reg soc_videooverlaysoc_core_ip_tx_target_unreachable = 1'd0;
wire [159:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header;
wire [15:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_value;
wire soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done;
reg [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r = 17'd0;
wire [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next0;
reg [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next0 = 17'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4checksum0 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next1;
reg [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next1 = 17'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4checksum1 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next2;
reg [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next2 = 17'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4checksum2 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next3;
reg [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next3 = 17'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4checksum3 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next4;
reg [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next4 = 17'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4checksum4 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next5;
reg [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next5 = 17'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4checksum5 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next6;
reg [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next6 = 17'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4checksum6 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next7;
reg [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next7 = 17'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4checksum7 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next8;
reg [16:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next8 = 17'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4checksum8 = 1'd0;
reg [3:0] soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_counter = 4'd0;
wire soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_counter_ce;
wire soc_videooverlaysoc_core_ip_tx_ce;
wire soc_videooverlaysoc_core_ip_tx_reset;
wire soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_valid;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_last;
wire [7:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_payload_data;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_payload_error = 1'd0;
wire [15:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_checksum;
wire [15:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_identification;
wire [3:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_ihl;
wire [7:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_protocol;
wire [31:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_sender_ip;
wire [31:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_target_ip;
wire [15:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_total_length;
wire [7:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_ttl;
wire [3:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_version;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid = 1'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_ready = 1'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_first = 1'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_last = 1'd0;
reg [15:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_ethernet_type = 16'd0;
reg [47:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_sender_mac = 48'd0;
reg [47:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_target_mac = 48'd0;
reg [7:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_last_be = 1'd0;
wire soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_error;
reg [159:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header = 160'd0;
reg [159:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header_reg = 160'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_load = 1'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_shift = 1'd0;
reg [4:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter = 5'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter_ce = 1'd0;
reg [7:0] soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer = 8'd0;
reg [47:0] soc_videooverlaysoc_core_ip_tx_target_mac = 48'd0;
wire soc_videooverlaysoc_core_ip_rx_sink_sink_valid;
wire soc_videooverlaysoc_core_ip_rx_sink_sink_ready;
wire soc_videooverlaysoc_core_ip_rx_sink_sink_first;
wire soc_videooverlaysoc_core_ip_rx_sink_sink_last;
wire [15:0] soc_videooverlaysoc_core_ip_rx_sink_sink_payload_ethernet_type;
wire [47:0] soc_videooverlaysoc_core_ip_rx_sink_sink_payload_sender_mac;
wire [47:0] soc_videooverlaysoc_core_ip_rx_sink_sink_payload_target_mac;
wire [7:0] soc_videooverlaysoc_core_ip_rx_sink_sink_payload_data;
wire soc_videooverlaysoc_core_ip_rx_sink_sink_payload_last_be;
wire soc_videooverlaysoc_core_ip_rx_sink_sink_payload_error;
reg soc_videooverlaysoc_core_ip_rx_source_source_valid = 1'd0;
wire soc_videooverlaysoc_core_ip_rx_source_source_ready;
reg soc_videooverlaysoc_core_ip_rx_source_source_first = 1'd0;
wire soc_videooverlaysoc_core_ip_rx_source_source_last;
wire [7:0] soc_videooverlaysoc_core_ip_rx_source_source_payload_data;
wire soc_videooverlaysoc_core_ip_rx_source_source_payload_error;
wire [15:0] soc_videooverlaysoc_core_ip_rx_source_source_param_length;
wire [7:0] soc_videooverlaysoc_core_ip_rx_source_source_param_protocol;
wire [31:0] soc_videooverlaysoc_core_ip_rx_source_source_param_ip_address;
wire soc_videooverlaysoc_core_ip_rx_depacketizer_sink_valid;
reg soc_videooverlaysoc_core_ip_rx_depacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_ip_rx_depacketizer_sink_first;
wire soc_videooverlaysoc_core_ip_rx_depacketizer_sink_last;
wire [15:0] soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_ethernet_type;
wire [47:0] soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_sender_mac;
wire [47:0] soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_target_mac;
wire [7:0] soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_data;
wire soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_last_be;
wire soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_error;
reg soc_videooverlaysoc_core_ip_rx_depacketizer_source_valid = 1'd0;
reg soc_videooverlaysoc_core_ip_rx_depacketizer_source_ready = 1'd0;
wire soc_videooverlaysoc_core_ip_rx_depacketizer_source_last;
wire [7:0] soc_videooverlaysoc_core_ip_rx_depacketizer_source_payload_data;
wire soc_videooverlaysoc_core_ip_rx_depacketizer_source_payload_error;
wire [15:0] soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_checksum;
wire [15:0] soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_identification;
wire [3:0] soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_ihl;
wire [7:0] soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_protocol;
wire [31:0] soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_sender_ip;
wire [31:0] soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_target_ip;
wire [15:0] soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_total_length;
wire [7:0] soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_ttl;
wire [3:0] soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_version;
wire [159:0] soc_videooverlaysoc_core_ip_rx_depacketizer_header;
reg [159:0] soc_videooverlaysoc_core_ip_rx_depacketizer_header_reg = 160'd0;
reg soc_videooverlaysoc_core_ip_rx_depacketizer_shift = 1'd0;
reg [4:0] soc_videooverlaysoc_core_ip_rx_depacketizer_counter = 5'd0;
reg soc_videooverlaysoc_core_ip_rx_depacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_ip_rx_depacketizer_counter_ce = 1'd0;
reg soc_videooverlaysoc_core_ip_rx_depacketizer_no_payload = 1'd0;
wire soc_videooverlaysoc_core_ip_rx_depacketizer_is_el;
wire [159:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header;
wire [15:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_value;
wire soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r = 17'd0;
wire [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next0;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next0 = 17'd0;
reg soc_videooverlaysoc_core_ip_rx_liteethipv4checksum0 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next1;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next1 = 17'd0;
reg soc_videooverlaysoc_core_ip_rx_liteethipv4checksum1 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next2;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next2 = 17'd0;
reg soc_videooverlaysoc_core_ip_rx_liteethipv4checksum2 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next3;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next3 = 17'd0;
reg soc_videooverlaysoc_core_ip_rx_liteethipv4checksum3 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next4;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next4 = 17'd0;
reg soc_videooverlaysoc_core_ip_rx_liteethipv4checksum4 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next5;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next5 = 17'd0;
reg soc_videooverlaysoc_core_ip_rx_liteethipv4checksum5 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next6;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next6 = 17'd0;
reg soc_videooverlaysoc_core_ip_rx_liteethipv4checksum6 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next7;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next7 = 17'd0;
reg soc_videooverlaysoc_core_ip_rx_liteethipv4checksum7 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next8;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next8 = 17'd0;
reg soc_videooverlaysoc_core_ip_rx_liteethipv4checksum8 = 1'd0;
wire [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next9;
reg [16:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next9 = 17'd0;
reg soc_videooverlaysoc_core_ip_rx_liteethipv4checksum9 = 1'd0;
reg [3:0] soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_counter = 4'd0;
wire soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_counter_ce;
wire soc_videooverlaysoc_core_ip_rx_ce;
wire soc_videooverlaysoc_core_ip_rx_reset;
reg soc_videooverlaysoc_core_ip_rx_valid = 1'd0;
wire soc_videooverlaysoc_core_ip_mac_port_sink_valid;
reg soc_videooverlaysoc_core_ip_mac_port_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_ip_mac_port_sink_first;
wire soc_videooverlaysoc_core_ip_mac_port_sink_last;
wire [15:0] soc_videooverlaysoc_core_ip_mac_port_sink_payload_ethernet_type;
wire [47:0] soc_videooverlaysoc_core_ip_mac_port_sink_payload_sender_mac;
wire [47:0] soc_videooverlaysoc_core_ip_mac_port_sink_payload_target_mac;
wire [7:0] soc_videooverlaysoc_core_ip_mac_port_sink_payload_data;
wire soc_videooverlaysoc_core_ip_mac_port_sink_payload_last_be;
wire soc_videooverlaysoc_core_ip_mac_port_sink_payload_error;
reg soc_videooverlaysoc_core_ip_mac_port_source_valid = 1'd0;
wire soc_videooverlaysoc_core_ip_mac_port_source_ready;
reg soc_videooverlaysoc_core_ip_mac_port_source_first = 1'd0;
reg soc_videooverlaysoc_core_ip_mac_port_source_last = 1'd0;
reg [15:0] soc_videooverlaysoc_core_ip_mac_port_source_payload_ethernet_type = 16'd0;
reg [47:0] soc_videooverlaysoc_core_ip_mac_port_source_payload_sender_mac = 48'd0;
reg [47:0] soc_videooverlaysoc_core_ip_mac_port_source_payload_target_mac = 48'd0;
reg [7:0] soc_videooverlaysoc_core_ip_mac_port_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_ip_mac_port_source_payload_last_be = 1'd0;
reg soc_videooverlaysoc_core_ip_mac_port_source_payload_error = 1'd0;
reg soc_videooverlaysoc_core_ip_crossbar_source_valid = 1'd0;
wire soc_videooverlaysoc_core_ip_crossbar_source_ready;
reg soc_videooverlaysoc_core_ip_crossbar_source_first = 1'd0;
reg soc_videooverlaysoc_core_ip_crossbar_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_ip_crossbar_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_ip_crossbar_source_payload_error = 1'd0;
reg [15:0] soc_videooverlaysoc_core_ip_crossbar_source_param_length = 16'd0;
reg [7:0] soc_videooverlaysoc_core_ip_crossbar_source_param_protocol = 8'd0;
reg [31:0] soc_videooverlaysoc_core_ip_crossbar_source_param_ip_address = 32'd0;
wire soc_videooverlaysoc_core_ip_crossbar_sink_valid;
reg soc_videooverlaysoc_core_ip_crossbar_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_ip_crossbar_sink_first;
wire soc_videooverlaysoc_core_ip_crossbar_sink_last;
wire [7:0] soc_videooverlaysoc_core_ip_crossbar_sink_payload_data;
wire soc_videooverlaysoc_core_ip_crossbar_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_ip_crossbar_sink_param_length;
wire [7:0] soc_videooverlaysoc_core_ip_crossbar_sink_param_protocol;
wire [31:0] soc_videooverlaysoc_core_ip_crossbar_sink_param_ip_address;
wire soc_videooverlaysoc_core_icmp_tx_sink_valid;
wire soc_videooverlaysoc_core_icmp_tx_sink_ready;
wire soc_videooverlaysoc_core_icmp_tx_sink_first;
wire soc_videooverlaysoc_core_icmp_tx_sink_last;
wire [7:0] soc_videooverlaysoc_core_icmp_tx_sink_payload_data;
wire soc_videooverlaysoc_core_icmp_tx_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_tx_sink_param_checksum;
wire [7:0] soc_videooverlaysoc_core_icmp_tx_sink_param_code;
wire [7:0] soc_videooverlaysoc_core_icmp_tx_sink_param_msgtype;
wire [31:0] soc_videooverlaysoc_core_icmp_tx_sink_param_quench;
wire [31:0] soc_videooverlaysoc_core_icmp_tx_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_icmp_tx_sink_param_length;
reg soc_videooverlaysoc_core_icmp_tx_source_valid = 1'd0;
wire soc_videooverlaysoc_core_icmp_tx_source_ready;
reg soc_videooverlaysoc_core_icmp_tx_source_first = 1'd0;
reg soc_videooverlaysoc_core_icmp_tx_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_icmp_tx_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_icmp_tx_source_payload_error = 1'd0;
reg [15:0] soc_videooverlaysoc_core_icmp_tx_source_param_length = 16'd0;
reg [7:0] soc_videooverlaysoc_core_icmp_tx_source_param_protocol = 8'd0;
reg [31:0] soc_videooverlaysoc_core_icmp_tx_source_param_ip_address = 32'd0;
wire soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_valid;
reg soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_last;
wire [7:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_payload_data;
reg soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_payload_error = 1'd0;
wire [15:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_checksum;
wire [7:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_code;
wire [7:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_msgtype;
wire [31:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_quench;
reg soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_valid = 1'd0;
reg soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_ready = 1'd0;
reg soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_first = 1'd0;
reg soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_payload_data = 8'd0;
wire soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_payload_error;
reg [15:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_param_length = 16'd0;
reg [7:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_param_protocol = 8'd0;
reg [31:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_param_ip_address = 32'd0;
reg [63:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header = 64'd0;
reg [63:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header_reg = 64'd0;
reg soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_load = 1'd0;
reg soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_shift = 1'd0;
reg [2:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter = 3'd0;
reg soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter_ce = 1'd0;
reg [7:0] soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer = 8'd0;
wire soc_videooverlaysoc_core_icmp_rx_sink_sink_valid;
wire soc_videooverlaysoc_core_icmp_rx_sink_sink_ready;
wire soc_videooverlaysoc_core_icmp_rx_sink_sink_first;
wire soc_videooverlaysoc_core_icmp_rx_sink_sink_last;
wire [7:0] soc_videooverlaysoc_core_icmp_rx_sink_sink_payload_data;
wire soc_videooverlaysoc_core_icmp_rx_sink_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_rx_sink_sink_param_length;
wire [7:0] soc_videooverlaysoc_core_icmp_rx_sink_sink_param_protocol;
wire [31:0] soc_videooverlaysoc_core_icmp_rx_sink_sink_param_ip_address;
reg soc_videooverlaysoc_core_icmp_rx_source_source_valid = 1'd0;
wire soc_videooverlaysoc_core_icmp_rx_source_source_ready;
reg soc_videooverlaysoc_core_icmp_rx_source_source_first = 1'd0;
wire soc_videooverlaysoc_core_icmp_rx_source_source_last;
wire [7:0] soc_videooverlaysoc_core_icmp_rx_source_source_payload_data;
wire soc_videooverlaysoc_core_icmp_rx_source_source_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_rx_source_source_param_checksum;
wire [7:0] soc_videooverlaysoc_core_icmp_rx_source_source_param_code;
wire [7:0] soc_videooverlaysoc_core_icmp_rx_source_source_param_msgtype;
wire [31:0] soc_videooverlaysoc_core_icmp_rx_source_source_param_quench;
wire [31:0] soc_videooverlaysoc_core_icmp_rx_source_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_icmp_rx_source_source_param_length;
wire soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_valid;
reg soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_first;
wire soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_last;
wire [7:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_payload_data;
wire soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_param_length;
wire [7:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_param_protocol;
wire [31:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_param_ip_address;
reg soc_videooverlaysoc_core_icmp_rx_depacketizer_source_valid = 1'd0;
reg soc_videooverlaysoc_core_icmp_rx_depacketizer_source_ready = 1'd0;
wire soc_videooverlaysoc_core_icmp_rx_depacketizer_source_last;
wire [7:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_source_payload_data;
wire soc_videooverlaysoc_core_icmp_rx_depacketizer_source_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_checksum;
wire [7:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_code;
wire [7:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_msgtype;
wire [31:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_quench;
wire [63:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_header;
reg [63:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_header_reg = 64'd0;
reg soc_videooverlaysoc_core_icmp_rx_depacketizer_shift = 1'd0;
reg [2:0] soc_videooverlaysoc_core_icmp_rx_depacketizer_counter = 3'd0;
reg soc_videooverlaysoc_core_icmp_rx_depacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_icmp_rx_depacketizer_counter_ce = 1'd0;
reg soc_videooverlaysoc_core_icmp_rx_depacketizer_no_payload = 1'd0;
wire soc_videooverlaysoc_core_icmp_rx_depacketizer_is_el;
reg soc_videooverlaysoc_core_icmp_rx_valid = 1'd0;
wire soc_videooverlaysoc_core_icmp_echo_sink_sink_valid;
wire soc_videooverlaysoc_core_icmp_echo_sink_sink_ready;
wire soc_videooverlaysoc_core_icmp_echo_sink_sink_first;
wire soc_videooverlaysoc_core_icmp_echo_sink_sink_last;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_sink_sink_payload_data;
wire soc_videooverlaysoc_core_icmp_echo_sink_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_sink_sink_param_checksum;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_sink_sink_param_code;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_sink_sink_param_msgtype;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_sink_sink_param_quench;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_sink_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_sink_sink_param_length;
wire soc_videooverlaysoc_core_icmp_echo_source_source_valid;
wire soc_videooverlaysoc_core_icmp_echo_source_source_ready;
wire soc_videooverlaysoc_core_icmp_echo_source_source_first;
wire soc_videooverlaysoc_core_icmp_echo_source_source_last;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_source_source_payload_data;
wire soc_videooverlaysoc_core_icmp_echo_source_source_payload_error;
reg [15:0] soc_videooverlaysoc_core_icmp_echo_source_source_param_checksum = 16'd0;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_source_source_param_code;
reg [7:0] soc_videooverlaysoc_core_icmp_echo_source_source_param_msgtype = 8'd0;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_source_source_param_quench;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_source_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_source_source_param_length;
wire soc_videooverlaysoc_core_icmp_echo_buffer_sink_valid;
wire soc_videooverlaysoc_core_icmp_echo_buffer_sink_ready;
wire soc_videooverlaysoc_core_icmp_echo_buffer_sink_first;
wire soc_videooverlaysoc_core_icmp_echo_buffer_sink_last;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_sink_payload_data;
wire soc_videooverlaysoc_core_icmp_echo_buffer_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_checksum;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_code;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_msgtype;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_quench;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_length;
wire soc_videooverlaysoc_core_icmp_echo_buffer_source_valid;
wire soc_videooverlaysoc_core_icmp_echo_buffer_source_ready;
wire soc_videooverlaysoc_core_icmp_echo_buffer_source_first;
wire soc_videooverlaysoc_core_icmp_echo_buffer_source_last;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_source_payload_data;
wire soc_videooverlaysoc_core_icmp_echo_buffer_source_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_buffer_source_param_checksum;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_source_param_code;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_source_param_msgtype;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_buffer_source_param_quench;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_buffer_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_buffer_source_param_length;
wire soc_videooverlaysoc_core_icmp_echo_buffer_re;
reg soc_videooverlaysoc_core_icmp_echo_buffer_readable = 1'd0;
wire soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_we;
wire soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_writable;
wire soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_re;
wire soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_readable;
wire [122:0] soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_din;
wire [122:0] soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_dout;
reg [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_level0 = 8'd0;
reg soc_videooverlaysoc_core_icmp_echo_buffer_replace = 1'd0;
reg [6:0] soc_videooverlaysoc_core_icmp_echo_buffer_produce = 7'd0;
reg [6:0] soc_videooverlaysoc_core_icmp_echo_buffer_consume = 7'd0;
reg [6:0] soc_videooverlaysoc_core_icmp_echo_buffer_wrport_adr = 7'd0;
wire [122:0] soc_videooverlaysoc_core_icmp_echo_buffer_wrport_dat_r;
wire soc_videooverlaysoc_core_icmp_echo_buffer_wrport_we;
wire [122:0] soc_videooverlaysoc_core_icmp_echo_buffer_wrport_dat_w;
wire soc_videooverlaysoc_core_icmp_echo_buffer_do_read;
wire [6:0] soc_videooverlaysoc_core_icmp_echo_buffer_rdport_adr;
wire [122:0] soc_videooverlaysoc_core_icmp_echo_buffer_rdport_dat_r;
wire soc_videooverlaysoc_core_icmp_echo_buffer_rdport_re;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_level1;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_payload_data;
wire soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_checksum;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_code;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_msgtype;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_quench;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_length;
wire soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_first;
wire soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_last;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_payload_data;
wire soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_checksum;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_code;
wire [7:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_msgtype;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_quench;
wire [31:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_length;
wire soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_first;
wire soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_last;
wire soc_videooverlaysoc_core_icmp_ip_port_sink_valid;
reg soc_videooverlaysoc_core_icmp_ip_port_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_icmp_ip_port_sink_first;
wire soc_videooverlaysoc_core_icmp_ip_port_sink_last;
wire [7:0] soc_videooverlaysoc_core_icmp_ip_port_sink_payload_data;
wire soc_videooverlaysoc_core_icmp_ip_port_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_icmp_ip_port_sink_param_length;
wire [7:0] soc_videooverlaysoc_core_icmp_ip_port_sink_param_protocol;
wire [31:0] soc_videooverlaysoc_core_icmp_ip_port_sink_param_ip_address;
reg soc_videooverlaysoc_core_icmp_ip_port_source_valid = 1'd0;
wire soc_videooverlaysoc_core_icmp_ip_port_source_ready;
reg soc_videooverlaysoc_core_icmp_ip_port_source_first = 1'd0;
reg soc_videooverlaysoc_core_icmp_ip_port_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_icmp_ip_port_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_icmp_ip_port_source_payload_error = 1'd0;
reg [15:0] soc_videooverlaysoc_core_icmp_ip_port_source_param_length = 16'd0;
reg [7:0] soc_videooverlaysoc_core_icmp_ip_port_source_param_protocol = 8'd0;
reg [31:0] soc_videooverlaysoc_core_icmp_ip_port_source_param_ip_address = 32'd0;
wire soc_videooverlaysoc_core_tx_sink_valid;
wire soc_videooverlaysoc_core_tx_sink_ready;
wire soc_videooverlaysoc_core_tx_sink_first;
wire soc_videooverlaysoc_core_tx_sink_last;
wire [7:0] soc_videooverlaysoc_core_tx_sink_payload_data;
wire soc_videooverlaysoc_core_tx_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_tx_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_core_tx_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_core_tx_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_tx_sink_param_length;
reg soc_videooverlaysoc_core_tx_source_valid = 1'd0;
wire soc_videooverlaysoc_core_tx_source_ready;
reg soc_videooverlaysoc_core_tx_source_first = 1'd0;
reg soc_videooverlaysoc_core_tx_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_tx_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_tx_source_payload_error = 1'd0;
reg [15:0] soc_videooverlaysoc_core_tx_source_param_length = 16'd0;
reg [7:0] soc_videooverlaysoc_core_tx_source_param_protocol = 8'd0;
reg [31:0] soc_videooverlaysoc_core_tx_source_param_ip_address = 32'd0;
wire soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_valid;
reg soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_last;
wire [7:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_payload_data;
reg soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_payload_error = 1'd0;
wire [15:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_checksum;
wire [15:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_dst_port;
wire [15:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_length;
wire [15:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_src_port;
reg soc_videooverlaysoc_core_tx_liteethudppacketizer_source_valid = 1'd0;
reg soc_videooverlaysoc_core_tx_liteethudppacketizer_source_ready = 1'd0;
reg soc_videooverlaysoc_core_tx_liteethudppacketizer_source_first = 1'd0;
reg soc_videooverlaysoc_core_tx_liteethudppacketizer_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_source_payload_data = 8'd0;
wire soc_videooverlaysoc_core_tx_liteethudppacketizer_source_payload_error;
reg [15:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_source_param_length = 16'd0;
reg [7:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_source_param_protocol = 8'd0;
reg [31:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_source_param_ip_address = 32'd0;
reg [63:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_header = 64'd0;
reg [63:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_header_reg = 64'd0;
reg soc_videooverlaysoc_core_tx_liteethudppacketizer_load = 1'd0;
reg soc_videooverlaysoc_core_tx_liteethudppacketizer_shift = 1'd0;
reg [2:0] soc_videooverlaysoc_core_tx_liteethudppacketizer_counter = 3'd0;
reg soc_videooverlaysoc_core_tx_liteethudppacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_tx_liteethudppacketizer_counter_ce = 1'd0;
reg [7:0] soc_videooverlaysoc_core_tx_liteethudppacketizer = 8'd0;
wire soc_videooverlaysoc_core_sink_sink_valid;
wire soc_videooverlaysoc_core_sink_sink_ready;
wire soc_videooverlaysoc_core_sink_sink_first;
wire soc_videooverlaysoc_core_sink_sink_last;
wire [7:0] soc_videooverlaysoc_core_sink_sink_payload_data;
wire soc_videooverlaysoc_core_sink_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_sink_sink_param_length;
wire [7:0] soc_videooverlaysoc_core_sink_sink_param_protocol;
wire [31:0] soc_videooverlaysoc_core_sink_sink_param_ip_address;
reg soc_videooverlaysoc_core_source_source_valid = 1'd0;
wire soc_videooverlaysoc_core_source_source_ready;
reg soc_videooverlaysoc_core_source_source_first = 1'd0;
wire soc_videooverlaysoc_core_source_source_last;
wire [7:0] soc_videooverlaysoc_core_source_source_payload_data;
wire soc_videooverlaysoc_core_source_source_payload_error;
wire [15:0] soc_videooverlaysoc_core_source_source_param_src_port;
wire [15:0] soc_videooverlaysoc_core_source_source_param_dst_port;
wire [31:0] soc_videooverlaysoc_core_source_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_source_source_param_length;
wire soc_videooverlaysoc_core_depacketizer_sink_valid;
reg soc_videooverlaysoc_core_depacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_depacketizer_sink_first;
wire soc_videooverlaysoc_core_depacketizer_sink_last;
wire [7:0] soc_videooverlaysoc_core_depacketizer_sink_payload_data;
wire soc_videooverlaysoc_core_depacketizer_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_depacketizer_sink_param_length;
wire [7:0] soc_videooverlaysoc_core_depacketizer_sink_param_protocol;
wire [31:0] soc_videooverlaysoc_core_depacketizer_sink_param_ip_address;
reg soc_videooverlaysoc_core_depacketizer_source_valid = 1'd0;
reg soc_videooverlaysoc_core_depacketizer_source_ready = 1'd0;
wire soc_videooverlaysoc_core_depacketizer_source_last;
wire [7:0] soc_videooverlaysoc_core_depacketizer_source_payload_data;
wire soc_videooverlaysoc_core_depacketizer_source_payload_error;
wire [15:0] soc_videooverlaysoc_core_depacketizer_source_param_checksum;
wire [15:0] soc_videooverlaysoc_core_depacketizer_source_param_dst_port;
wire [15:0] soc_videooverlaysoc_core_depacketizer_source_param_length;
wire [15:0] soc_videooverlaysoc_core_depacketizer_source_param_src_port;
wire [63:0] soc_videooverlaysoc_core_depacketizer_header;
reg [63:0] soc_videooverlaysoc_core_depacketizer_header_reg = 64'd0;
reg soc_videooverlaysoc_core_depacketizer_shift = 1'd0;
reg [2:0] soc_videooverlaysoc_core_depacketizer_counter = 3'd0;
reg soc_videooverlaysoc_core_depacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_core_depacketizer_counter_ce = 1'd0;
reg soc_videooverlaysoc_core_depacketizer_no_payload = 1'd0;
wire soc_videooverlaysoc_core_depacketizer_is_el;
reg soc_videooverlaysoc_core_valid = 1'd0;
wire soc_videooverlaysoc_core_ip_port_sink_valid;
reg soc_videooverlaysoc_core_ip_port_sink_ready = 1'd0;
wire soc_videooverlaysoc_core_ip_port_sink_first;
wire soc_videooverlaysoc_core_ip_port_sink_last;
wire [7:0] soc_videooverlaysoc_core_ip_port_sink_payload_data;
wire soc_videooverlaysoc_core_ip_port_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_ip_port_sink_param_length;
wire [7:0] soc_videooverlaysoc_core_ip_port_sink_param_protocol;
wire [31:0] soc_videooverlaysoc_core_ip_port_sink_param_ip_address;
reg soc_videooverlaysoc_core_ip_port_source_valid = 1'd0;
wire soc_videooverlaysoc_core_ip_port_source_ready;
reg soc_videooverlaysoc_core_ip_port_source_first = 1'd0;
reg soc_videooverlaysoc_core_ip_port_source_last = 1'd0;
reg [7:0] soc_videooverlaysoc_core_ip_port_source_payload_data = 8'd0;
reg soc_videooverlaysoc_core_ip_port_source_payload_error = 1'd0;
reg [15:0] soc_videooverlaysoc_core_ip_port_source_param_length = 16'd0;
reg [7:0] soc_videooverlaysoc_core_ip_port_source_param_protocol = 8'd0;
reg [31:0] soc_videooverlaysoc_core_ip_port_source_param_ip_address = 32'd0;
wire soc_videooverlaysoc_core_crossbar_source_valid;
wire soc_videooverlaysoc_core_crossbar_source_ready;
wire soc_videooverlaysoc_core_crossbar_source_first;
wire soc_videooverlaysoc_core_crossbar_source_last;
wire [7:0] soc_videooverlaysoc_core_crossbar_source_payload_data;
wire soc_videooverlaysoc_core_crossbar_source_payload_error;
wire [15:0] soc_videooverlaysoc_core_crossbar_source_param_src_port;
wire [15:0] soc_videooverlaysoc_core_crossbar_source_param_dst_port;
wire [31:0] soc_videooverlaysoc_core_crossbar_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_crossbar_source_param_length;
wire soc_videooverlaysoc_core_crossbar_sink_valid;
wire soc_videooverlaysoc_core_crossbar_sink_ready;
wire soc_videooverlaysoc_core_crossbar_sink_first;
wire soc_videooverlaysoc_core_crossbar_sink_last;
wire [7:0] soc_videooverlaysoc_core_crossbar_sink_payload_data;
wire soc_videooverlaysoc_core_crossbar_sink_payload_error;
wire [15:0] soc_videooverlaysoc_core_crossbar_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_core_crossbar_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_core_crossbar_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_core_crossbar_sink_param_length;
wire etherbone_clk;
wire etherbone_rst;
reg soc_videooverlaysoc_packet_sink_valid = 1'd0;
wire soc_videooverlaysoc_packet_sink_ready;
reg soc_videooverlaysoc_packet_sink_first = 1'd0;
reg soc_videooverlaysoc_packet_sink_last = 1'd0;
reg [31:0] soc_videooverlaysoc_packet_sink_payload_data = 32'd0;
reg [3:0] soc_videooverlaysoc_packet_sink_payload_error = 4'd0;
reg [3:0] soc_videooverlaysoc_packet_sink_param_addr_size = 4'd0;
reg soc_videooverlaysoc_packet_sink_param_nr = 1'd0;
reg soc_videooverlaysoc_packet_sink_param_pf = 1'd0;
reg [3:0] soc_videooverlaysoc_packet_sink_param_port_size = 4'd0;
reg soc_videooverlaysoc_packet_sink_param_pr = 1'd0;
reg [15:0] soc_videooverlaysoc_packet_sink_param_src_port = 16'd0;
reg [15:0] soc_videooverlaysoc_packet_sink_param_dst_port = 16'd0;
reg [31:0] soc_videooverlaysoc_packet_sink_param_ip_address = 32'd0;
reg [15:0] soc_videooverlaysoc_packet_sink_param_length = 16'd0;
reg soc_videooverlaysoc_packet_source_valid = 1'd0;
wire soc_videooverlaysoc_packet_source_ready;
reg soc_videooverlaysoc_packet_source_first = 1'd0;
reg soc_videooverlaysoc_packet_source_last = 1'd0;
reg [31:0] soc_videooverlaysoc_packet_source_payload_data = 32'd0;
reg [3:0] soc_videooverlaysoc_packet_source_payload_error = 4'd0;
reg [15:0] soc_videooverlaysoc_packet_source_param_src_port = 16'd0;
reg [15:0] soc_videooverlaysoc_packet_source_param_dst_port = 16'd0;
reg [31:0] soc_videooverlaysoc_packet_source_param_ip_address = 32'd0;
reg [15:0] soc_videooverlaysoc_packet_source_param_length = 16'd0;
wire soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_valid;
reg soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_last;
wire [31:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_payload_data;
reg [3:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_payload_error = 4'd0;
wire [3:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_addr_size;
wire [15:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_magic;
wire soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_nr;
wire soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_pf;
wire [3:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_port_size;
wire soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_pr;
wire [3:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_version;
reg soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_valid = 1'd0;
reg soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_ready = 1'd0;
reg soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_first = 1'd0;
reg soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_last = 1'd0;
reg [31:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_payload_data = 32'd0;
wire [3:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_payload_error;
reg [15:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_param_src_port = 16'd0;
reg [15:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_param_dst_port = 16'd0;
reg [31:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_param_ip_address = 32'd0;
reg [15:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_param_length = 16'd0;
reg [63:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header = 64'd0;
reg [63:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header_reg = 64'd0;
reg soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_load = 1'd0;
reg soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_shift = 1'd0;
reg soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter = 1'd0;
reg soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter_ce = 1'd0;
reg [31:0] soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer = 32'd0;
wire soc_videooverlaysoc_packet_sink_sink_valid;
wire soc_videooverlaysoc_packet_sink_sink_ready;
wire soc_videooverlaysoc_packet_sink_sink_first;
wire soc_videooverlaysoc_packet_sink_sink_last;
wire [31:0] soc_videooverlaysoc_packet_sink_sink_payload_data;
wire [3:0] soc_videooverlaysoc_packet_sink_sink_payload_error;
wire [15:0] soc_videooverlaysoc_packet_sink_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_sink_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_sink_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_sink_sink_param_length;
reg soc_videooverlaysoc_packet_source_source_valid = 1'd0;
reg soc_videooverlaysoc_packet_source_source_ready = 1'd0;
reg soc_videooverlaysoc_packet_source_source_first = 1'd0;
wire soc_videooverlaysoc_packet_source_source_last;
wire [31:0] soc_videooverlaysoc_packet_source_source_payload_data;
reg [3:0] soc_videooverlaysoc_packet_source_source_payload_error = 4'd0;
reg [3:0] soc_videooverlaysoc_packet_source_source_param_addr_size = 4'd0;
wire soc_videooverlaysoc_packet_source_source_param_nr;
wire soc_videooverlaysoc_packet_source_source_param_pf;
reg [3:0] soc_videooverlaysoc_packet_source_source_param_port_size = 4'd0;
wire soc_videooverlaysoc_packet_source_source_param_pr;
wire [15:0] soc_videooverlaysoc_packet_source_source_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_source_source_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_source_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_source_source_param_length;
wire soc_videooverlaysoc_packet_depacketizer_sink_valid;
reg soc_videooverlaysoc_packet_depacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_packet_depacketizer_sink_first;
wire soc_videooverlaysoc_packet_depacketizer_sink_last;
wire [31:0] soc_videooverlaysoc_packet_depacketizer_sink_payload_data;
wire [3:0] soc_videooverlaysoc_packet_depacketizer_sink_payload_error;
wire [15:0] soc_videooverlaysoc_packet_depacketizer_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_depacketizer_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_depacketizer_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_depacketizer_sink_param_length;
reg soc_videooverlaysoc_packet_depacketizer_source_valid = 1'd0;
reg soc_videooverlaysoc_packet_depacketizer_source_ready = 1'd0;
wire soc_videooverlaysoc_packet_depacketizer_source_last;
wire [31:0] soc_videooverlaysoc_packet_depacketizer_source_payload_data;
wire [3:0] soc_videooverlaysoc_packet_depacketizer_source_payload_error;
wire [3:0] soc_videooverlaysoc_packet_depacketizer_source_param_addr_size;
wire [15:0] soc_videooverlaysoc_packet_depacketizer_source_param_magic;
wire soc_videooverlaysoc_packet_depacketizer_source_param_nr;
wire soc_videooverlaysoc_packet_depacketizer_source_param_pf;
wire [3:0] soc_videooverlaysoc_packet_depacketizer_source_param_port_size;
wire soc_videooverlaysoc_packet_depacketizer_source_param_pr;
wire [3:0] soc_videooverlaysoc_packet_depacketizer_source_param_version;
wire [63:0] soc_videooverlaysoc_packet_depacketizer_header;
reg [63:0] soc_videooverlaysoc_packet_depacketizer_header_reg = 64'd0;
reg soc_videooverlaysoc_packet_depacketizer_shift = 1'd0;
reg soc_videooverlaysoc_packet_depacketizer_counter = 1'd0;
reg soc_videooverlaysoc_packet_depacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_packet_depacketizer_counter_ce = 1'd0;
reg soc_videooverlaysoc_packet_depacketizer_no_payload = 1'd0;
wire soc_videooverlaysoc_packet_depacketizer_is_el;
reg soc_videooverlaysoc_packet_valid = 1'd0;
wire soc_videooverlaysoc_packet_user_port_sink_valid;
wire soc_videooverlaysoc_packet_user_port_sink_ready;
wire soc_videooverlaysoc_packet_user_port_sink_first;
wire soc_videooverlaysoc_packet_user_port_sink_last;
wire [31:0] soc_videooverlaysoc_packet_user_port_sink_payload_data;
wire [3:0] soc_videooverlaysoc_packet_user_port_sink_payload_error;
wire [15:0] soc_videooverlaysoc_packet_user_port_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_user_port_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_user_port_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_user_port_sink_param_length;
wire soc_videooverlaysoc_packet_user_port_source_valid;
wire soc_videooverlaysoc_packet_user_port_source_ready;
wire soc_videooverlaysoc_packet_user_port_source_first;
wire soc_videooverlaysoc_packet_user_port_source_last;
wire [31:0] soc_videooverlaysoc_packet_user_port_source_payload_data;
wire [3:0] soc_videooverlaysoc_packet_user_port_source_payload_error;
wire [15:0] soc_videooverlaysoc_packet_user_port_source_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_user_port_source_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_user_port_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_user_port_source_param_length;
wire soc_videooverlaysoc_packet_internal_port_sink_valid;
wire soc_videooverlaysoc_packet_internal_port_sink_ready;
wire soc_videooverlaysoc_packet_internal_port_sink_first;
wire soc_videooverlaysoc_packet_internal_port_sink_last;
wire [7:0] soc_videooverlaysoc_packet_internal_port_sink_payload_data;
wire soc_videooverlaysoc_packet_internal_port_sink_payload_error;
wire [15:0] soc_videooverlaysoc_packet_internal_port_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_internal_port_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_internal_port_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_internal_port_sink_param_length;
wire soc_videooverlaysoc_packet_internal_port_source_valid;
wire soc_videooverlaysoc_packet_internal_port_source_ready;
wire soc_videooverlaysoc_packet_internal_port_source_first;
wire soc_videooverlaysoc_packet_internal_port_source_last;
wire [7:0] soc_videooverlaysoc_packet_internal_port_source_payload_data;
wire soc_videooverlaysoc_packet_internal_port_source_payload_error;
wire [15:0] soc_videooverlaysoc_packet_internal_port_source_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_internal_port_source_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_internal_port_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_internal_port_source_param_length;
wire soc_videooverlaysoc_packet_tx_cdc_sink_valid;
wire soc_videooverlaysoc_packet_tx_cdc_sink_ready;
wire soc_videooverlaysoc_packet_tx_cdc_sink_first;
wire soc_videooverlaysoc_packet_tx_cdc_sink_last;
wire [31:0] soc_videooverlaysoc_packet_tx_cdc_sink_payload_data;
wire [3:0] soc_videooverlaysoc_packet_tx_cdc_sink_payload_error;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_tx_cdc_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_sink_param_length;
wire soc_videooverlaysoc_packet_tx_cdc_source_valid;
wire soc_videooverlaysoc_packet_tx_cdc_source_ready;
wire soc_videooverlaysoc_packet_tx_cdc_source_first;
wire soc_videooverlaysoc_packet_tx_cdc_source_last;
wire [31:0] soc_videooverlaysoc_packet_tx_cdc_source_payload_data;
wire [3:0] soc_videooverlaysoc_packet_tx_cdc_source_payload_error;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_source_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_source_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_tx_cdc_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_source_param_length;
wire soc_videooverlaysoc_packet_tx_cdc_asyncfifo_we;
wire soc_videooverlaysoc_packet_tx_cdc_asyncfifo_writable;
wire soc_videooverlaysoc_packet_tx_cdc_asyncfifo_re;
wire soc_videooverlaysoc_packet_tx_cdc_asyncfifo_readable;
wire [117:0] soc_videooverlaysoc_packet_tx_cdc_asyncfifo_din;
wire [117:0] soc_videooverlaysoc_packet_tx_cdc_asyncfifo_dout;
wire soc_videooverlaysoc_packet_tx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [2:0] soc_videooverlaysoc_packet_tx_cdc_graycounter0_q = 3'd0;
wire [2:0] soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_next;
reg [2:0] soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_binary = 3'd0;
reg [2:0] soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_next_binary = 3'd0;
wire soc_videooverlaysoc_packet_tx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [2:0] soc_videooverlaysoc_packet_tx_cdc_graycounter1_q = 3'd0;
wire [2:0] soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next;
reg [2:0] soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_binary = 3'd0;
reg [2:0] soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next_binary = 3'd0;
wire [2:0] soc_videooverlaysoc_packet_tx_cdc_produce_rdomain;
wire [2:0] soc_videooverlaysoc_packet_tx_cdc_consume_wdomain;
wire [1:0] soc_videooverlaysoc_packet_tx_cdc_wrport_adr;
wire [117:0] soc_videooverlaysoc_packet_tx_cdc_wrport_dat_r;
wire soc_videooverlaysoc_packet_tx_cdc_wrport_we;
wire [117:0] soc_videooverlaysoc_packet_tx_cdc_wrport_dat_w;
wire [1:0] soc_videooverlaysoc_packet_tx_cdc_rdport_adr;
wire [117:0] soc_videooverlaysoc_packet_tx_cdc_rdport_dat_r;
wire [31:0] soc_videooverlaysoc_packet_tx_cdc_fifo_in_payload_data;
wire [3:0] soc_videooverlaysoc_packet_tx_cdc_fifo_in_payload_error;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_length;
wire soc_videooverlaysoc_packet_tx_cdc_fifo_in_first;
wire soc_videooverlaysoc_packet_tx_cdc_fifo_in_last;
wire [31:0] soc_videooverlaysoc_packet_tx_cdc_fifo_out_payload_data;
wire [3:0] soc_videooverlaysoc_packet_tx_cdc_fifo_out_payload_error;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_length;
wire soc_videooverlaysoc_packet_tx_cdc_fifo_out_first;
wire soc_videooverlaysoc_packet_tx_cdc_fifo_out_last;
wire soc_videooverlaysoc_packet_tx_converter_sink_valid;
wire soc_videooverlaysoc_packet_tx_converter_sink_ready;
wire soc_videooverlaysoc_packet_tx_converter_sink_first;
wire soc_videooverlaysoc_packet_tx_converter_sink_last;
wire [31:0] soc_videooverlaysoc_packet_tx_converter_sink_payload_data;
wire [3:0] soc_videooverlaysoc_packet_tx_converter_sink_payload_error;
wire [15:0] soc_videooverlaysoc_packet_tx_converter_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_tx_converter_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_tx_converter_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_tx_converter_sink_param_length;
wire soc_videooverlaysoc_packet_tx_converter_source_valid;
wire soc_videooverlaysoc_packet_tx_converter_source_ready;
wire soc_videooverlaysoc_packet_tx_converter_source_first;
wire soc_videooverlaysoc_packet_tx_converter_source_last;
wire [7:0] soc_videooverlaysoc_packet_tx_converter_source_payload_data;
wire soc_videooverlaysoc_packet_tx_converter_source_payload_error;
wire [15:0] soc_videooverlaysoc_packet_tx_converter_source_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_tx_converter_source_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_tx_converter_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_tx_converter_source_param_length;
wire soc_videooverlaysoc_packet_tx_converter_converter_sink_valid;
wire soc_videooverlaysoc_packet_tx_converter_converter_sink_ready;
wire soc_videooverlaysoc_packet_tx_converter_converter_sink_first;
wire soc_videooverlaysoc_packet_tx_converter_converter_sink_last;
reg [35:0] soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data = 36'd0;
wire soc_videooverlaysoc_packet_tx_converter_converter_source_valid;
wire soc_videooverlaysoc_packet_tx_converter_converter_source_ready;
wire soc_videooverlaysoc_packet_tx_converter_converter_source_first;
wire soc_videooverlaysoc_packet_tx_converter_converter_source_last;
reg [8:0] soc_videooverlaysoc_packet_tx_converter_converter_source_payload_data = 9'd0;
wire soc_videooverlaysoc_packet_tx_converter_converter_source_payload_valid_token_count;
reg [1:0] soc_videooverlaysoc_packet_tx_converter_converter_mux = 2'd0;
wire soc_videooverlaysoc_packet_tx_converter_converter_first;
wire soc_videooverlaysoc_packet_tx_converter_converter_last;
wire soc_videooverlaysoc_packet_tx_converter_source_source_valid;
wire soc_videooverlaysoc_packet_tx_converter_source_source_ready;
wire soc_videooverlaysoc_packet_tx_converter_source_source_first;
wire soc_videooverlaysoc_packet_tx_converter_source_source_last;
wire [8:0] soc_videooverlaysoc_packet_tx_converter_source_source_payload_data;
wire soc_videooverlaysoc_packet_rx_converter_sink_valid;
wire soc_videooverlaysoc_packet_rx_converter_sink_ready;
wire soc_videooverlaysoc_packet_rx_converter_sink_first;
wire soc_videooverlaysoc_packet_rx_converter_sink_last;
wire [7:0] soc_videooverlaysoc_packet_rx_converter_sink_payload_data;
wire soc_videooverlaysoc_packet_rx_converter_sink_payload_error;
wire [15:0] soc_videooverlaysoc_packet_rx_converter_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_rx_converter_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_rx_converter_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_rx_converter_sink_param_length;
wire soc_videooverlaysoc_packet_rx_converter_source_valid;
wire soc_videooverlaysoc_packet_rx_converter_source_ready;
wire soc_videooverlaysoc_packet_rx_converter_source_first;
wire soc_videooverlaysoc_packet_rx_converter_source_last;
reg [31:0] soc_videooverlaysoc_packet_rx_converter_source_payload_data = 32'd0;
reg [3:0] soc_videooverlaysoc_packet_rx_converter_source_payload_error = 4'd0;
reg [15:0] soc_videooverlaysoc_packet_rx_converter_source_param_src_port = 16'd0;
reg [15:0] soc_videooverlaysoc_packet_rx_converter_source_param_dst_port = 16'd0;
reg [31:0] soc_videooverlaysoc_packet_rx_converter_source_param_ip_address = 32'd0;
reg [15:0] soc_videooverlaysoc_packet_rx_converter_source_param_length = 16'd0;
wire soc_videooverlaysoc_packet_rx_converter_converter_sink_valid;
wire soc_videooverlaysoc_packet_rx_converter_converter_sink_ready;
wire soc_videooverlaysoc_packet_rx_converter_converter_sink_first;
wire soc_videooverlaysoc_packet_rx_converter_converter_sink_last;
wire [8:0] soc_videooverlaysoc_packet_rx_converter_converter_sink_payload_data;
wire soc_videooverlaysoc_packet_rx_converter_converter_source_valid;
wire soc_videooverlaysoc_packet_rx_converter_converter_source_ready;
reg soc_videooverlaysoc_packet_rx_converter_converter_source_first = 1'd0;
reg soc_videooverlaysoc_packet_rx_converter_converter_source_last = 1'd0;
reg [35:0] soc_videooverlaysoc_packet_rx_converter_converter_source_payload_data = 36'd0;
reg [2:0] soc_videooverlaysoc_packet_rx_converter_converter_source_payload_valid_token_count = 3'd0;
reg [1:0] soc_videooverlaysoc_packet_rx_converter_converter_demux = 2'd0;
wire soc_videooverlaysoc_packet_rx_converter_converter_load_part;
reg soc_videooverlaysoc_packet_rx_converter_converter_strobe_all = 1'd0;
wire soc_videooverlaysoc_packet_rx_converter_source_source_valid;
wire soc_videooverlaysoc_packet_rx_converter_source_source_ready;
wire soc_videooverlaysoc_packet_rx_converter_source_source_first;
wire soc_videooverlaysoc_packet_rx_converter_source_source_last;
wire [35:0] soc_videooverlaysoc_packet_rx_converter_source_source_payload_data;
wire soc_videooverlaysoc_packet_rx_cdc_sink_valid;
wire soc_videooverlaysoc_packet_rx_cdc_sink_ready;
wire soc_videooverlaysoc_packet_rx_cdc_sink_first;
wire soc_videooverlaysoc_packet_rx_cdc_sink_last;
wire [31:0] soc_videooverlaysoc_packet_rx_cdc_sink_payload_data;
wire [3:0] soc_videooverlaysoc_packet_rx_cdc_sink_payload_error;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_rx_cdc_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_sink_param_length;
wire soc_videooverlaysoc_packet_rx_cdc_source_valid;
wire soc_videooverlaysoc_packet_rx_cdc_source_ready;
wire soc_videooverlaysoc_packet_rx_cdc_source_first;
wire soc_videooverlaysoc_packet_rx_cdc_source_last;
wire [31:0] soc_videooverlaysoc_packet_rx_cdc_source_payload_data;
wire [3:0] soc_videooverlaysoc_packet_rx_cdc_source_payload_error;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_source_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_source_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_rx_cdc_source_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_source_param_length;
wire soc_videooverlaysoc_packet_rx_cdc_asyncfifo_we;
wire soc_videooverlaysoc_packet_rx_cdc_asyncfifo_writable;
wire soc_videooverlaysoc_packet_rx_cdc_asyncfifo_re;
wire soc_videooverlaysoc_packet_rx_cdc_asyncfifo_readable;
wire [117:0] soc_videooverlaysoc_packet_rx_cdc_asyncfifo_din;
wire [117:0] soc_videooverlaysoc_packet_rx_cdc_asyncfifo_dout;
wire soc_videooverlaysoc_packet_rx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [2:0] soc_videooverlaysoc_packet_rx_cdc_graycounter0_q = 3'd0;
wire [2:0] soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_next;
reg [2:0] soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_binary = 3'd0;
reg [2:0] soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_next_binary = 3'd0;
wire soc_videooverlaysoc_packet_rx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [2:0] soc_videooverlaysoc_packet_rx_cdc_graycounter1_q = 3'd0;
wire [2:0] soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next;
reg [2:0] soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_binary = 3'd0;
reg [2:0] soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next_binary = 3'd0;
wire [2:0] soc_videooverlaysoc_packet_rx_cdc_produce_rdomain;
wire [2:0] soc_videooverlaysoc_packet_rx_cdc_consume_wdomain;
wire [1:0] soc_videooverlaysoc_packet_rx_cdc_wrport_adr;
wire [117:0] soc_videooverlaysoc_packet_rx_cdc_wrport_dat_r;
wire soc_videooverlaysoc_packet_rx_cdc_wrport_we;
wire [117:0] soc_videooverlaysoc_packet_rx_cdc_wrport_dat_w;
wire [1:0] soc_videooverlaysoc_packet_rx_cdc_rdport_adr;
wire [117:0] soc_videooverlaysoc_packet_rx_cdc_rdport_dat_r;
wire [31:0] soc_videooverlaysoc_packet_rx_cdc_fifo_in_payload_data;
wire [3:0] soc_videooverlaysoc_packet_rx_cdc_fifo_in_payload_error;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_length;
wire soc_videooverlaysoc_packet_rx_cdc_fifo_in_first;
wire soc_videooverlaysoc_packet_rx_cdc_fifo_in_last;
wire [31:0] soc_videooverlaysoc_packet_rx_cdc_fifo_out_payload_data;
wire [3:0] soc_videooverlaysoc_packet_rx_cdc_fifo_out_payload_error;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_src_port;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_dst_port;
wire [31:0] soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_ip_address;
wire [15:0] soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_length;
wire soc_videooverlaysoc_packet_rx_cdc_fifo_out_first;
wire soc_videooverlaysoc_packet_rx_cdc_fifo_out_last;
reg soc_videooverlaysoc_probe_sink_valid = 1'd0;
reg soc_videooverlaysoc_probe_sink_ready = 1'd0;
reg soc_videooverlaysoc_probe_sink_first = 1'd0;
reg soc_videooverlaysoc_probe_sink_last = 1'd0;
reg [31:0] soc_videooverlaysoc_probe_sink_payload_data = 32'd0;
reg [3:0] soc_videooverlaysoc_probe_sink_payload_error = 4'd0;
reg [3:0] soc_videooverlaysoc_probe_sink_param_addr_size = 4'd0;
reg soc_videooverlaysoc_probe_sink_param_nr = 1'd0;
reg soc_videooverlaysoc_probe_sink_param_pf = 1'd0;
reg [3:0] soc_videooverlaysoc_probe_sink_param_port_size = 4'd0;
reg soc_videooverlaysoc_probe_sink_param_pr = 1'd0;
reg [15:0] soc_videooverlaysoc_probe_sink_param_src_port = 16'd0;
reg [15:0] soc_videooverlaysoc_probe_sink_param_dst_port = 16'd0;
reg [31:0] soc_videooverlaysoc_probe_sink_param_ip_address = 32'd0;
reg [15:0] soc_videooverlaysoc_probe_sink_param_length = 16'd0;
reg soc_videooverlaysoc_probe_source_valid = 1'd0;
reg soc_videooverlaysoc_probe_source_ready = 1'd0;
reg soc_videooverlaysoc_probe_source_first = 1'd0;
reg soc_videooverlaysoc_probe_source_last = 1'd0;
reg [31:0] soc_videooverlaysoc_probe_source_payload_data = 32'd0;
reg [3:0] soc_videooverlaysoc_probe_source_payload_error = 4'd0;
reg [3:0] soc_videooverlaysoc_probe_source_param_addr_size = 4'd0;
reg soc_videooverlaysoc_probe_source_param_nr = 1'd0;
reg soc_videooverlaysoc_probe_source_param_pf = 1'd0;
reg [3:0] soc_videooverlaysoc_probe_source_param_port_size = 4'd0;
reg soc_videooverlaysoc_probe_source_param_pr = 1'd0;
reg [15:0] soc_videooverlaysoc_probe_source_param_src_port = 16'd0;
reg [15:0] soc_videooverlaysoc_probe_source_param_dst_port = 16'd0;
reg [31:0] soc_videooverlaysoc_probe_source_param_ip_address = 32'd0;
reg [15:0] soc_videooverlaysoc_probe_source_param_length = 16'd0;
reg soc_videooverlaysoc_record_sink_sink_valid = 1'd0;
wire soc_videooverlaysoc_record_sink_sink_ready;
reg soc_videooverlaysoc_record_sink_sink_first = 1'd0;
reg soc_videooverlaysoc_record_sink_sink_last = 1'd0;
reg [31:0] soc_videooverlaysoc_record_sink_sink_payload_data = 32'd0;
reg [3:0] soc_videooverlaysoc_record_sink_sink_payload_error = 4'd0;
reg [3:0] soc_videooverlaysoc_record_sink_sink_param_addr_size = 4'd0;
reg soc_videooverlaysoc_record_sink_sink_param_nr = 1'd0;
reg soc_videooverlaysoc_record_sink_sink_param_pf = 1'd0;
reg [3:0] soc_videooverlaysoc_record_sink_sink_param_port_size = 4'd0;
reg soc_videooverlaysoc_record_sink_sink_param_pr = 1'd0;
reg [15:0] soc_videooverlaysoc_record_sink_sink_param_src_port = 16'd0;
reg [15:0] soc_videooverlaysoc_record_sink_sink_param_dst_port = 16'd0;
reg [31:0] soc_videooverlaysoc_record_sink_sink_param_ip_address = 32'd0;
reg [15:0] soc_videooverlaysoc_record_sink_sink_param_length = 16'd0;
wire soc_videooverlaysoc_record_source_source_valid;
reg soc_videooverlaysoc_record_source_source_ready = 1'd0;
wire soc_videooverlaysoc_record_source_source_first;
wire soc_videooverlaysoc_record_source_source_last;
wire [31:0] soc_videooverlaysoc_record_source_source_payload_data;
wire [3:0] soc_videooverlaysoc_record_source_source_payload_error;
wire [3:0] soc_videooverlaysoc_record_source_source_param_addr_size;
wire soc_videooverlaysoc_record_source_source_param_nr;
wire soc_videooverlaysoc_record_source_source_param_pf;
wire [3:0] soc_videooverlaysoc_record_source_source_param_port_size;
wire soc_videooverlaysoc_record_source_source_param_pr;
wire [15:0] soc_videooverlaysoc_record_source_source_param_src_port;
wire [15:0] soc_videooverlaysoc_record_source_source_param_dst_port;
reg [31:0] soc_videooverlaysoc_record_source_source_param_ip_address = 32'd0;
reg [15:0] soc_videooverlaysoc_record_source_source_param_length = 16'd0;
wire soc_videooverlaysoc_record_depacketizer_sink_valid;
reg soc_videooverlaysoc_record_depacketizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_record_depacketizer_sink_first;
wire soc_videooverlaysoc_record_depacketizer_sink_last;
wire [31:0] soc_videooverlaysoc_record_depacketizer_sink_payload_data;
wire [3:0] soc_videooverlaysoc_record_depacketizer_sink_payload_error;
wire [3:0] soc_videooverlaysoc_record_depacketizer_sink_param_addr_size;
wire soc_videooverlaysoc_record_depacketizer_sink_param_nr;
wire soc_videooverlaysoc_record_depacketizer_sink_param_pf;
wire [3:0] soc_videooverlaysoc_record_depacketizer_sink_param_port_size;
wire soc_videooverlaysoc_record_depacketizer_sink_param_pr;
wire [15:0] soc_videooverlaysoc_record_depacketizer_sink_param_src_port;
wire [15:0] soc_videooverlaysoc_record_depacketizer_sink_param_dst_port;
wire [31:0] soc_videooverlaysoc_record_depacketizer_sink_param_ip_address;
wire [15:0] soc_videooverlaysoc_record_depacketizer_sink_param_length;
reg soc_videooverlaysoc_record_depacketizer_source_valid = 1'd0;
wire soc_videooverlaysoc_record_depacketizer_source_ready;
reg soc_videooverlaysoc_record_depacketizer_source_first = 1'd0;
wire soc_videooverlaysoc_record_depacketizer_source_last;
wire [31:0] soc_videooverlaysoc_record_depacketizer_source_payload_data;
wire [3:0] soc_videooverlaysoc_record_depacketizer_source_payload_error;
wire soc_videooverlaysoc_record_depacketizer_source_param_bca;
wire [7:0] soc_videooverlaysoc_record_depacketizer_source_param_byte_enable;
wire soc_videooverlaysoc_record_depacketizer_source_param_cyc;
wire soc_videooverlaysoc_record_depacketizer_source_param_rca;
wire [7:0] soc_videooverlaysoc_record_depacketizer_source_param_rcount;
wire soc_videooverlaysoc_record_depacketizer_source_param_rff;
wire soc_videooverlaysoc_record_depacketizer_source_param_wca;
wire [7:0] soc_videooverlaysoc_record_depacketizer_source_param_wcount;
wire soc_videooverlaysoc_record_depacketizer_source_param_wff;
wire [31:0] soc_videooverlaysoc_record_depacketizer_header;
reg [31:0] soc_videooverlaysoc_record_depacketizer_header_reg = 32'd0;
reg soc_videooverlaysoc_record_depacketizer_shift = 1'd0;
reg soc_videooverlaysoc_record_depacketizer_counter = 1'd0;
reg soc_videooverlaysoc_record_depacketizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_record_depacketizer_counter_ce = 1'd0;
reg soc_videooverlaysoc_record_depacketizer_no_payload = 1'd0;
wire soc_videooverlaysoc_record_depacketizer_is_el;
wire soc_videooverlaysoc_record_receiver_sink_sink_valid;
wire soc_videooverlaysoc_record_receiver_sink_sink_ready;
wire soc_videooverlaysoc_record_receiver_sink_sink_first;
wire soc_videooverlaysoc_record_receiver_sink_sink_last;
reg [31:0] soc_videooverlaysoc_record_receiver_sink_sink_payload_data = 32'd0;
wire [3:0] soc_videooverlaysoc_record_receiver_sink_sink_payload_error;
wire soc_videooverlaysoc_record_receiver_sink_sink_param_bca;
wire [7:0] soc_videooverlaysoc_record_receiver_sink_sink_param_byte_enable;
wire soc_videooverlaysoc_record_receiver_sink_sink_param_cyc;
wire soc_videooverlaysoc_record_receiver_sink_sink_param_rca;
wire [7:0] soc_videooverlaysoc_record_receiver_sink_sink_param_rcount;
wire soc_videooverlaysoc_record_receiver_sink_sink_param_rff;
wire soc_videooverlaysoc_record_receiver_sink_sink_param_wca;
wire [7:0] soc_videooverlaysoc_record_receiver_sink_sink_param_wcount;
wire soc_videooverlaysoc_record_receiver_sink_sink_param_wff;
reg soc_videooverlaysoc_record_receiver_source_source_valid = 1'd0;
wire soc_videooverlaysoc_record_receiver_source_source_ready;
reg soc_videooverlaysoc_record_receiver_source_source_first = 1'd0;
reg soc_videooverlaysoc_record_receiver_source_source_last = 1'd0;
reg [31:0] soc_videooverlaysoc_record_receiver_source_source_payload_addr = 32'd0;
reg [31:0] soc_videooverlaysoc_record_receiver_source_source_payload_data = 32'd0;
reg soc_videooverlaysoc_record_receiver_source_source_param_we = 1'd0;
reg [7:0] soc_videooverlaysoc_record_receiver_source_source_param_count = 8'd0;
reg [31:0] soc_videooverlaysoc_record_receiver_source_source_param_base_addr = 32'd0;
reg [3:0] soc_videooverlaysoc_record_receiver_source_source_param_be = 4'd0;
wire soc_videooverlaysoc_record_receiver_fifo_sink_valid;
wire soc_videooverlaysoc_record_receiver_fifo_sink_ready;
wire soc_videooverlaysoc_record_receiver_fifo_sink_first;
wire soc_videooverlaysoc_record_receiver_fifo_sink_last;
wire [31:0] soc_videooverlaysoc_record_receiver_fifo_sink_payload_data;
wire [3:0] soc_videooverlaysoc_record_receiver_fifo_sink_payload_error;
wire soc_videooverlaysoc_record_receiver_fifo_sink_param_bca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_sink_param_byte_enable;
wire soc_videooverlaysoc_record_receiver_fifo_sink_param_cyc;
wire soc_videooverlaysoc_record_receiver_fifo_sink_param_rca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_sink_param_rcount;
wire soc_videooverlaysoc_record_receiver_fifo_sink_param_rff;
wire soc_videooverlaysoc_record_receiver_fifo_sink_param_wca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_sink_param_wcount;
wire soc_videooverlaysoc_record_receiver_fifo_sink_param_wff;
wire soc_videooverlaysoc_record_receiver_fifo_source_valid;
reg soc_videooverlaysoc_record_receiver_fifo_source_ready = 1'd0;
wire soc_videooverlaysoc_record_receiver_fifo_source_first;
wire soc_videooverlaysoc_record_receiver_fifo_source_last;
wire [31:0] soc_videooverlaysoc_record_receiver_fifo_source_payload_data;
wire [3:0] soc_videooverlaysoc_record_receiver_fifo_source_payload_error;
wire soc_videooverlaysoc_record_receiver_fifo_source_param_bca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_source_param_byte_enable;
wire soc_videooverlaysoc_record_receiver_fifo_source_param_cyc;
wire soc_videooverlaysoc_record_receiver_fifo_source_param_rca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_source_param_rcount;
wire soc_videooverlaysoc_record_receiver_fifo_source_param_rff;
wire soc_videooverlaysoc_record_receiver_fifo_source_param_wca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_source_param_wcount;
wire soc_videooverlaysoc_record_receiver_fifo_source_param_wff;
wire soc_videooverlaysoc_record_receiver_fifo_re;
reg soc_videooverlaysoc_record_receiver_fifo_readable = 1'd0;
wire soc_videooverlaysoc_record_receiver_fifo_syncfifo_we;
wire soc_videooverlaysoc_record_receiver_fifo_syncfifo_writable;
wire soc_videooverlaysoc_record_receiver_fifo_syncfifo_re;
wire soc_videooverlaysoc_record_receiver_fifo_syncfifo_readable;
wire [67:0] soc_videooverlaysoc_record_receiver_fifo_syncfifo_din;
wire [67:0] soc_videooverlaysoc_record_receiver_fifo_syncfifo_dout;
reg [2:0] soc_videooverlaysoc_record_receiver_fifo_level0 = 3'd0;
reg soc_videooverlaysoc_record_receiver_fifo_replace = 1'd0;
reg [1:0] soc_videooverlaysoc_record_receiver_fifo_produce = 2'd0;
reg [1:0] soc_videooverlaysoc_record_receiver_fifo_consume = 2'd0;
reg [1:0] soc_videooverlaysoc_record_receiver_fifo_wrport_adr = 2'd0;
wire [67:0] soc_videooverlaysoc_record_receiver_fifo_wrport_dat_r;
wire soc_videooverlaysoc_record_receiver_fifo_wrport_we;
wire [67:0] soc_videooverlaysoc_record_receiver_fifo_wrport_dat_w;
wire soc_videooverlaysoc_record_receiver_fifo_do_read;
wire [1:0] soc_videooverlaysoc_record_receiver_fifo_rdport_adr;
wire [67:0] soc_videooverlaysoc_record_receiver_fifo_rdport_dat_r;
wire soc_videooverlaysoc_record_receiver_fifo_rdport_re;
wire [2:0] soc_videooverlaysoc_record_receiver_fifo_level1;
wire [31:0] soc_videooverlaysoc_record_receiver_fifo_fifo_in_payload_data;
wire [3:0] soc_videooverlaysoc_record_receiver_fifo_fifo_in_payload_error;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_bca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_byte_enable;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_cyc;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_rca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_rcount;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_rff;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_wca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_wcount;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_wff;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_in_first;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_in_last;
wire [31:0] soc_videooverlaysoc_record_receiver_fifo_fifo_out_payload_data;
wire [3:0] soc_videooverlaysoc_record_receiver_fifo_fifo_out_payload_error;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_bca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_byte_enable;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_cyc;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_rca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_rcount;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_rff;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_wca;
wire [7:0] soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_wcount;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_wff;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_out_first;
wire soc_videooverlaysoc_record_receiver_fifo_fifo_out_last;
reg [31:0] soc_videooverlaysoc_record_receiver_base_addr = 32'd0;
reg soc_videooverlaysoc_record_receiver_base_addr_update = 1'd0;
reg [8:0] soc_videooverlaysoc_record_receiver_counter = 9'd0;
reg soc_videooverlaysoc_record_receiver_counter_reset = 1'd0;
reg soc_videooverlaysoc_record_receiver_counter_ce = 1'd0;
reg soc_videooverlaysoc_record_first = 1'd1;
reg [31:0] soc_videooverlaysoc_record_last_ip_address = 32'd0;
wire soc_videooverlaysoc_record_sender_sink_sink_valid;
wire soc_videooverlaysoc_record_sender_sink_sink_ready;
wire soc_videooverlaysoc_record_sender_sink_sink_first;
wire soc_videooverlaysoc_record_sender_sink_sink_last;
wire [31:0] soc_videooverlaysoc_record_sender_sink_sink_payload_addr;
wire [31:0] soc_videooverlaysoc_record_sender_sink_sink_payload_data;
wire soc_videooverlaysoc_record_sender_sink_sink_param_we;
wire [7:0] soc_videooverlaysoc_record_sender_sink_sink_param_count;
wire [31:0] soc_videooverlaysoc_record_sender_sink_sink_param_base_addr;
wire [3:0] soc_videooverlaysoc_record_sender_sink_sink_param_be;
reg soc_videooverlaysoc_record_sender_source_source_valid = 1'd0;
wire soc_videooverlaysoc_record_sender_source_source_ready;
reg soc_videooverlaysoc_record_sender_source_source_first = 1'd0;
reg soc_videooverlaysoc_record_sender_source_source_last = 1'd0;
reg [31:0] soc_videooverlaysoc_record_sender_source_source_payload_data = 32'd0;
reg [3:0] soc_videooverlaysoc_record_sender_source_source_payload_error = 4'd0;
reg soc_videooverlaysoc_record_sender_source_source_param_bca = 1'd0;
reg [7:0] soc_videooverlaysoc_record_sender_source_source_param_byte_enable = 8'd0;
reg soc_videooverlaysoc_record_sender_source_source_param_cyc = 1'd0;
reg soc_videooverlaysoc_record_sender_source_source_param_rca = 1'd0;
reg [7:0] soc_videooverlaysoc_record_sender_source_source_param_rcount = 8'd0;
reg soc_videooverlaysoc_record_sender_source_source_param_rff = 1'd0;
reg soc_videooverlaysoc_record_sender_source_source_param_wca = 1'd0;
reg [7:0] soc_videooverlaysoc_record_sender_source_source_param_wcount = 8'd0;
reg soc_videooverlaysoc_record_sender_source_source_param_wff = 1'd0;
wire soc_videooverlaysoc_record_sender_fifo_sink_valid;
wire soc_videooverlaysoc_record_sender_fifo_sink_ready;
wire soc_videooverlaysoc_record_sender_fifo_sink_first;
wire soc_videooverlaysoc_record_sender_fifo_sink_last;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_sink_payload_addr;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_sink_payload_data;
wire soc_videooverlaysoc_record_sender_fifo_sink_param_we;
wire [7:0] soc_videooverlaysoc_record_sender_fifo_sink_param_count;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_sink_param_base_addr;
wire [3:0] soc_videooverlaysoc_record_sender_fifo_sink_param_be;
wire soc_videooverlaysoc_record_sender_fifo_source_valid;
reg soc_videooverlaysoc_record_sender_fifo_source_ready = 1'd0;
wire soc_videooverlaysoc_record_sender_fifo_source_first;
wire soc_videooverlaysoc_record_sender_fifo_source_last;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_source_payload_addr;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_source_payload_data;
wire soc_videooverlaysoc_record_sender_fifo_source_param_we;
wire [7:0] soc_videooverlaysoc_record_sender_fifo_source_param_count;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_source_param_base_addr;
wire [3:0] soc_videooverlaysoc_record_sender_fifo_source_param_be;
wire soc_videooverlaysoc_record_sender_fifo_re;
reg soc_videooverlaysoc_record_sender_fifo_readable = 1'd0;
wire soc_videooverlaysoc_record_sender_fifo_syncfifo_we;
wire soc_videooverlaysoc_record_sender_fifo_syncfifo_writable;
wire soc_videooverlaysoc_record_sender_fifo_syncfifo_re;
wire soc_videooverlaysoc_record_sender_fifo_syncfifo_readable;
wire [110:0] soc_videooverlaysoc_record_sender_fifo_syncfifo_din;
wire [110:0] soc_videooverlaysoc_record_sender_fifo_syncfifo_dout;
reg [2:0] soc_videooverlaysoc_record_sender_fifo_level0 = 3'd0;
reg soc_videooverlaysoc_record_sender_fifo_replace = 1'd0;
reg [1:0] soc_videooverlaysoc_record_sender_fifo_produce = 2'd0;
reg [1:0] soc_videooverlaysoc_record_sender_fifo_consume = 2'd0;
reg [1:0] soc_videooverlaysoc_record_sender_fifo_wrport_adr = 2'd0;
wire [110:0] soc_videooverlaysoc_record_sender_fifo_wrport_dat_r;
wire soc_videooverlaysoc_record_sender_fifo_wrport_we;
wire [110:0] soc_videooverlaysoc_record_sender_fifo_wrport_dat_w;
wire soc_videooverlaysoc_record_sender_fifo_do_read;
wire [1:0] soc_videooverlaysoc_record_sender_fifo_rdport_adr;
wire [110:0] soc_videooverlaysoc_record_sender_fifo_rdport_dat_r;
wire soc_videooverlaysoc_record_sender_fifo_rdport_re;
wire [2:0] soc_videooverlaysoc_record_sender_fifo_level1;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_fifo_in_payload_addr;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_fifo_in_payload_data;
wire soc_videooverlaysoc_record_sender_fifo_fifo_in_param_we;
wire [7:0] soc_videooverlaysoc_record_sender_fifo_fifo_in_param_count;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_fifo_in_param_base_addr;
wire [3:0] soc_videooverlaysoc_record_sender_fifo_fifo_in_param_be;
wire soc_videooverlaysoc_record_sender_fifo_fifo_in_first;
wire soc_videooverlaysoc_record_sender_fifo_fifo_in_last;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_fifo_out_payload_addr;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_fifo_out_payload_data;
wire soc_videooverlaysoc_record_sender_fifo_fifo_out_param_we;
wire [7:0] soc_videooverlaysoc_record_sender_fifo_fifo_out_param_count;
wire [31:0] soc_videooverlaysoc_record_sender_fifo_fifo_out_param_base_addr;
wire [3:0] soc_videooverlaysoc_record_sender_fifo_fifo_out_param_be;
wire soc_videooverlaysoc_record_sender_fifo_fifo_out_first;
wire soc_videooverlaysoc_record_sender_fifo_fifo_out_last;
reg soc_videooverlaysoc_record_sender_data_sel = 1'd0;
wire soc_videooverlaysoc_record_packetizer_sink_valid;
reg soc_videooverlaysoc_record_packetizer_sink_ready = 1'd0;
wire soc_videooverlaysoc_record_packetizer_sink_first;
wire soc_videooverlaysoc_record_packetizer_sink_last;
reg [31:0] soc_videooverlaysoc_record_packetizer_sink_payload_data = 32'd0;
wire [3:0] soc_videooverlaysoc_record_packetizer_sink_payload_error;
wire soc_videooverlaysoc_record_packetizer_sink_param_bca;
wire [7:0] soc_videooverlaysoc_record_packetizer_sink_param_byte_enable;
wire soc_videooverlaysoc_record_packetizer_sink_param_cyc;
wire soc_videooverlaysoc_record_packetizer_sink_param_rca;
wire [7:0] soc_videooverlaysoc_record_packetizer_sink_param_rcount;
wire soc_videooverlaysoc_record_packetizer_sink_param_rff;
wire soc_videooverlaysoc_record_packetizer_sink_param_wca;
wire [7:0] soc_videooverlaysoc_record_packetizer_sink_param_wcount;
wire soc_videooverlaysoc_record_packetizer_sink_param_wff;
reg soc_videooverlaysoc_record_packetizer_source_valid = 1'd0;
wire soc_videooverlaysoc_record_packetizer_source_ready;
reg soc_videooverlaysoc_record_packetizer_source_first = 1'd0;
reg soc_videooverlaysoc_record_packetizer_source_last = 1'd0;
reg [31:0] soc_videooverlaysoc_record_packetizer_source_payload_data = 32'd0;
wire [3:0] soc_videooverlaysoc_record_packetizer_source_payload_error;
reg [3:0] soc_videooverlaysoc_record_packetizer_source_param_addr_size = 4'd0;
reg soc_videooverlaysoc_record_packetizer_source_param_nr = 1'd0;
reg soc_videooverlaysoc_record_packetizer_source_param_pf = 1'd0;
reg [3:0] soc_videooverlaysoc_record_packetizer_source_param_port_size = 4'd0;
reg soc_videooverlaysoc_record_packetizer_source_param_pr = 1'd0;
reg [15:0] soc_videooverlaysoc_record_packetizer_source_param_src_port = 16'd0;
reg [15:0] soc_videooverlaysoc_record_packetizer_source_param_dst_port = 16'd0;
reg [31:0] soc_videooverlaysoc_record_packetizer_source_param_ip_address = 32'd0;
reg [15:0] soc_videooverlaysoc_record_packetizer_source_param_length = 16'd0;
reg [31:0] soc_videooverlaysoc_record_packetizer_header = 32'd0;
reg [31:0] soc_videooverlaysoc_record_packetizer_header_reg = 32'd0;
reg soc_videooverlaysoc_record_packetizer_load = 1'd0;
reg soc_videooverlaysoc_record_packetizer_counter = 1'd0;
reg soc_videooverlaysoc_record_packetizer_counter_reset = 1'd0;
reg soc_videooverlaysoc_record_packetizer_counter_ce = 1'd0;
wire soc_videooverlaysoc_dispatcher_sel0;
reg soc_videooverlaysoc_dispatcher_first = 1'd1;
reg soc_videooverlaysoc_dispatcher_last = 1'd0;
wire soc_videooverlaysoc_dispatcher_ongoing0;
reg soc_videooverlaysoc_dispatcher_ongoing1 = 1'd0;
reg soc_videooverlaysoc_dispatcher_sel1 = 1'd0;
reg soc_videooverlaysoc_dispatcher_sel_ongoing = 1'd0;
reg [1:0] soc_videooverlaysoc_request = 2'd0;
reg soc_videooverlaysoc_grant = 1'd0;
reg soc_videooverlaysoc_status0_first = 1'd1;
reg soc_videooverlaysoc_status0_last = 1'd0;
wire soc_videooverlaysoc_status0_ongoing0;
reg soc_videooverlaysoc_status0_ongoing1 = 1'd0;
reg soc_videooverlaysoc_status1_first = 1'd1;
reg soc_videooverlaysoc_status1_last = 1'd0;
wire soc_videooverlaysoc_status1_ongoing0;
reg soc_videooverlaysoc_status1_ongoing1 = 1'd0;
wire soc_videooverlaysoc_wishbone_sink_valid;
reg soc_videooverlaysoc_wishbone_sink_ready = 1'd0;
wire soc_videooverlaysoc_wishbone_sink_first;
wire soc_videooverlaysoc_wishbone_sink_last;
wire [31:0] soc_videooverlaysoc_wishbone_sink_payload_addr;
wire [31:0] soc_videooverlaysoc_wishbone_sink_payload_data;
wire soc_videooverlaysoc_wishbone_sink_param_we;
wire [7:0] soc_videooverlaysoc_wishbone_sink_param_count;
wire [31:0] soc_videooverlaysoc_wishbone_sink_param_base_addr;
wire [3:0] soc_videooverlaysoc_wishbone_sink_param_be;
reg soc_videooverlaysoc_wishbone_source_valid = 1'd0;
wire soc_videooverlaysoc_wishbone_source_ready;
reg soc_videooverlaysoc_wishbone_source_first = 1'd0;
reg soc_videooverlaysoc_wishbone_source_last = 1'd0;
reg [31:0] soc_videooverlaysoc_wishbone_source_payload_addr = 32'd0;
reg [31:0] soc_videooverlaysoc_wishbone_source_payload_data = 32'd0;
reg soc_videooverlaysoc_wishbone_source_param_we = 1'd0;
reg [7:0] soc_videooverlaysoc_wishbone_source_param_count = 8'd0;
reg [31:0] soc_videooverlaysoc_wishbone_source_param_base_addr = 32'd0;
reg [3:0] soc_videooverlaysoc_wishbone_source_param_be = 4'd0;
reg [29:0] soc_videooverlaysoc_wishbone_bus_adr = 30'd0;
reg [31:0] soc_videooverlaysoc_wishbone_bus_dat_w = 32'd0;
wire [31:0] soc_videooverlaysoc_wishbone_bus_dat_r;
reg [3:0] soc_videooverlaysoc_wishbone_bus_sel = 4'd0;
reg soc_videooverlaysoc_wishbone_bus_cyc = 1'd0;
reg soc_videooverlaysoc_wishbone_bus_stb = 1'd0;
wire soc_videooverlaysoc_wishbone_bus_ack;
reg soc_videooverlaysoc_wishbone_bus_we = 1'd0;
reg [2:0] soc_videooverlaysoc_wishbone_bus_cti = 3'd0;
reg [1:0] soc_videooverlaysoc_wishbone_bus_bte = 2'd0;
wire soc_videooverlaysoc_wishbone_bus_err;
reg soc_videooverlaysoc_wishbone_data_update = 1'd0;
reg [1:0] vns_refresher_state = 2'd0;
reg [1:0] vns_refresher_next_state = 2'd0;
reg [3:0] vns_bankmachine0_state = 4'd0;
reg [3:0] vns_bankmachine0_next_state = 4'd0;
reg [3:0] vns_bankmachine1_state = 4'd0;
reg [3:0] vns_bankmachine1_next_state = 4'd0;
reg [3:0] vns_bankmachine2_state = 4'd0;
reg [3:0] vns_bankmachine2_next_state = 4'd0;
reg [3:0] vns_bankmachine3_state = 4'd0;
reg [3:0] vns_bankmachine3_next_state = 4'd0;
reg [3:0] vns_bankmachine4_state = 4'd0;
reg [3:0] vns_bankmachine4_next_state = 4'd0;
reg [3:0] vns_bankmachine5_state = 4'd0;
reg [3:0] vns_bankmachine5_next_state = 4'd0;
reg [3:0] vns_bankmachine6_state = 4'd0;
reg [3:0] vns_bankmachine6_next_state = 4'd0;
reg [3:0] vns_bankmachine7_state = 4'd0;
reg [3:0] vns_bankmachine7_next_state = 4'd0;
reg [3:0] vns_multiplexer_state = 4'd0;
reg [3:0] vns_multiplexer_next_state = 4'd0;
wire [2:0] vns_roundrobin0_request;
reg [1:0] vns_roundrobin0_grant = 2'd0;
wire vns_roundrobin0_ce;
wire [2:0] vns_roundrobin1_request;
reg [1:0] vns_roundrobin1_grant = 2'd0;
wire vns_roundrobin1_ce;
wire [2:0] vns_roundrobin2_request;
reg [1:0] vns_roundrobin2_grant = 2'd0;
wire vns_roundrobin2_ce;
wire [2:0] vns_roundrobin3_request;
reg [1:0] vns_roundrobin3_grant = 2'd0;
wire vns_roundrobin3_ce;
wire [2:0] vns_roundrobin4_request;
reg [1:0] vns_roundrobin4_grant = 2'd0;
wire vns_roundrobin4_ce;
wire [2:0] vns_roundrobin5_request;
reg [1:0] vns_roundrobin5_grant = 2'd0;
wire vns_roundrobin5_ce;
wire [2:0] vns_roundrobin6_request;
reg [1:0] vns_roundrobin6_grant = 2'd0;
wire vns_roundrobin6_ce;
wire [2:0] vns_roundrobin7_request;
reg [1:0] vns_roundrobin7_grant = 2'd0;
wire vns_roundrobin7_ce;
reg [2:0] vns_rbank = 3'd0;
reg [2:0] vns_wbank = 3'd0;
reg vns_locked0 = 1'd0;
reg vns_locked1 = 1'd0;
reg vns_locked2 = 1'd0;
reg vns_locked3 = 1'd0;
reg vns_locked4 = 1'd0;
reg vns_locked5 = 1'd0;
reg vns_locked6 = 1'd0;
reg vns_locked7 = 1'd0;
reg vns_locked8 = 1'd0;
reg vns_locked9 = 1'd0;
reg vns_locked10 = 1'd0;
reg vns_locked11 = 1'd0;
reg vns_locked12 = 1'd0;
reg vns_locked13 = 1'd0;
reg vns_locked14 = 1'd0;
reg vns_locked15 = 1'd0;
reg vns_locked16 = 1'd0;
reg vns_locked17 = 1'd0;
reg vns_locked18 = 1'd0;
reg vns_locked19 = 1'd0;
reg vns_locked20 = 1'd0;
reg vns_locked21 = 1'd0;
reg vns_locked22 = 1'd0;
reg vns_locked23 = 1'd0;
reg vns_new_master_wdata_ready0 = 1'd0;
reg vns_new_master_wdata_ready1 = 1'd0;
reg vns_new_master_wdata_ready2 = 1'd0;
reg vns_new_master_wdata_ready3 = 1'd0;
reg vns_new_master_wdata_ready4 = 1'd0;
reg vns_new_master_wdata_ready5 = 1'd0;
reg vns_new_master_wdata_ready6 = 1'd0;
reg vns_new_master_wdata_ready7 = 1'd0;
reg vns_new_master_wdata_ready8 = 1'd0;
reg vns_new_master_rdata_valid0 = 1'd0;
reg vns_new_master_rdata_valid1 = 1'd0;
reg vns_new_master_rdata_valid2 = 1'd0;
reg vns_new_master_rdata_valid3 = 1'd0;
reg vns_new_master_rdata_valid4 = 1'd0;
reg vns_new_master_rdata_valid5 = 1'd0;
reg vns_new_master_rdata_valid6 = 1'd0;
reg vns_new_master_rdata_valid7 = 1'd0;
reg vns_new_master_rdata_valid8 = 1'd0;
reg vns_new_master_rdata_valid9 = 1'd0;
reg vns_new_master_rdata_valid10 = 1'd0;
reg vns_new_master_rdata_valid11 = 1'd0;
reg vns_new_master_rdata_valid12 = 1'd0;
reg vns_new_master_rdata_valid13 = 1'd0;
reg vns_new_master_rdata_valid14 = 1'd0;
reg vns_new_master_rdata_valid15 = 1'd0;
reg vns_new_master_rdata_valid16 = 1'd0;
reg vns_new_master_rdata_valid17 = 1'd0;
reg vns_new_master_rdata_valid18 = 1'd0;
reg vns_new_master_rdata_valid19 = 1'd0;
reg vns_new_master_rdata_valid20 = 1'd0;
reg vns_new_master_rdata_valid21 = 1'd0;
reg vns_new_master_rdata_valid22 = 1'd0;
reg vns_new_master_rdata_valid23 = 1'd0;
reg vns_new_master_rdata_valid24 = 1'd0;
reg vns_new_master_rdata_valid25 = 1'd0;
reg vns_new_master_rdata_valid26 = 1'd0;
reg vns_new_master_rdata_valid27 = 1'd0;
reg vns_new_master_rdata_valid28 = 1'd0;
reg vns_new_master_rdata_valid29 = 1'd0;
reg [2:0] vns_fullmemorywe_state = 3'd0;
reg [2:0] vns_fullmemorywe_next_state = 3'd0;
reg [1:0] vns_litedramwishbone2native_state = 2'd0;
reg [1:0] vns_litedramwishbone2native_next_state = 2'd0;
reg [3:0] vns_edid0_state = 4'd0;
reg [3:0] vns_edid0_next_state = 4'd0;
reg [2:0] vns_clockdomainsrenamer0_state0 = 3'd0;
reg [2:0] vns_clockdomainsrenamer0_next_state0 = 3'd0;
reg [3:0] vns_edid1_state = 4'd0;
reg [3:0] vns_edid1_next_state = 4'd0;
reg [2:0] vns_clockdomainsrenamer1_state0 = 3'd0;
reg [2:0] vns_clockdomainsrenamer1_next_state0 = 3'd0;
reg [1:0] vns_dma_state = 2'd0;
reg [1:0] vns_dma_next_state = 2'd0;
reg [1:0] vns_videooutcore_state = 2'd0;
reg [1:0] vns_videooutcore_next_state = 2'd0;
reg [26:0] soc_videooverlaysoc_hdmi_core_out0_dmareader_offset_next_value = 27'd0;
reg soc_videooverlaysoc_hdmi_core_out0_dmareader_offset_next_value_ce = 1'd0;
reg vns_clockdomainsrenamer0_state1 = 1'd0;
reg vns_clockdomainsrenamer0_next_state1 = 1'd0;
reg vns_clockdomainsrenamer1_liteethmac_liteethmacgap_state = 1'd0;
reg vns_clockdomainsrenamer1_liteethmac_liteethmacgap_next_state = 1'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_next_state = 2'd0;
reg vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_state = 1'd0;
reg vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_next_state = 1'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_next_state = 2'd0;
reg vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_state = 1'd0;
reg vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_next_state = 1'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_request = 2'd0;
reg vns_clockdomainsrenamer1_liteethmac_grant = 1'd0;
reg vns_clockdomainsrenamer1_liteethmac_status0_first = 1'd1;
reg vns_clockdomainsrenamer1_liteethmac_status0_last = 1'd0;
wire vns_clockdomainsrenamer1_liteethmac_status0_ongoing0;
reg vns_clockdomainsrenamer1_liteethmac_status0_ongoing1 = 1'd0;
reg vns_clockdomainsrenamer1_liteethmac_status1_first = 1'd1;
reg vns_clockdomainsrenamer1_liteethmac_status1_last = 1'd0;
wire vns_clockdomainsrenamer1_liteethmac_status1_ongoing0;
reg vns_clockdomainsrenamer1_liteethmac_status1_ongoing1 = 1'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_sel0 = 2'd0;
reg vns_clockdomainsrenamer1_liteethmac_first = 1'd1;
reg vns_clockdomainsrenamer1_liteethmac_last = 1'd0;
wire vns_clockdomainsrenamer1_liteethmac_ongoing0;
reg vns_clockdomainsrenamer1_liteethmac_ongoing1 = 1'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_sel1 = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_sel_ongoing = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_next_state = 2'd0;
reg vns_clockdomainsrenamer1_liteetharptx_fsm_state = 1'd0;
reg vns_clockdomainsrenamer1_liteetharptx_fsm_next_state = 1'd0;
reg [1:0] vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteetharprx_fsm_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteetharprx_fsm_next_state = 2'd0;
reg [2:0] vns_clockdomainsrenamer1_state1 = 3'd0;
reg [2:0] vns_clockdomainsrenamer1_next_state1 = 3'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_next_state = 2'd0;
reg [2:0] vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_state = 3'd0;
reg [2:0] vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_next_state = 3'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethip_request = 2'd0;
reg vns_clockdomainsrenamer1_liteethip_grant = 1'd0;
reg vns_clockdomainsrenamer1_liteethip_status0_first = 1'd1;
reg vns_clockdomainsrenamer1_liteethip_status0_last = 1'd0;
wire vns_clockdomainsrenamer1_liteethip_status0_ongoing0;
reg vns_clockdomainsrenamer1_liteethip_status0_ongoing1 = 1'd0;
reg vns_clockdomainsrenamer1_liteethip_status1_first = 1'd1;
reg vns_clockdomainsrenamer1_liteethip_status1_last = 1'd0;
wire vns_clockdomainsrenamer1_liteethip_status1_ongoing0;
reg vns_clockdomainsrenamer1_liteethip_status1_ongoing1 = 1'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethip_sel0 = 2'd0;
reg vns_clockdomainsrenamer1_liteethip_first = 1'd1;
reg vns_clockdomainsrenamer1_liteethip_last = 1'd0;
wire vns_clockdomainsrenamer1_liteethip_ongoing0;
reg vns_clockdomainsrenamer1_liteethip_ongoing1 = 1'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethip_sel1 = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethip_sel_ongoing = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_next_state = 2'd0;
reg vns_clockdomainsrenamer1_liteethicmptx_fsm_state = 1'd0;
reg vns_clockdomainsrenamer1_liteethicmptx_fsm_next_state = 1'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethicmprx_fsm_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethicmprx_fsm_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_next_state = 2'd0;
reg vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_state = 1'd0;
reg vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_next_state = 1'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_next_state = 2'd0;
reg vns_clockdomainsrenamer1_liteethudp_sel = 1'd0;
reg [1:0] vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_state = 2'd0;
reg [1:0] vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_next_state = 2'd0;
reg vns_liteethetherbonepackettx_fsm_state = 1'd0;
reg vns_liteethetherbonepackettx_fsm_next_state = 1'd0;
reg [1:0] vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_state = 2'd0;
reg [1:0] vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_next_state = 2'd0;
reg [1:0] vns_liteethetherbonepacketrx_fsm_state = 2'd0;
reg [1:0] vns_liteethetherbonepacketrx_fsm_next_state = 2'd0;
reg vns_liteethetherboneprobe_state = 1'd0;
reg vns_liteethetherboneprobe_next_state = 1'd0;
reg vns_liteethetherbonerecorddepacketizer_state = 1'd0;
reg vns_liteethetherbonerecorddepacketizer_next_state = 1'd0;
reg [1:0] vns_liteethetherbonerecordreceiver_state = 2'd0;
reg [1:0] vns_liteethetherbonerecordreceiver_next_state = 2'd0;
reg [1:0] vns_liteethetherbonerecordsender_state = 2'd0;
reg [1:0] vns_liteethetherbonerecordsender_next_state = 2'd0;
reg vns_liteethetherbonerecordpacketizer_state = 1'd0;
reg vns_liteethetherbonerecordpacketizer_next_state = 1'd0;
reg [1:0] vns_liteethetherbonewishbonemaster_state = 2'd0;
reg [1:0] vns_liteethetherbonewishbonemaster_next_state = 2'd0;
wire vns_wb_sdram_con_request;
wire vns_wb_sdram_con_grant;
wire [29:0] vns_videooverlaysoc_shared_adr;
wire [31:0] vns_videooverlaysoc_shared_dat_w;
reg [31:0] vns_videooverlaysoc_shared_dat_r = 32'd0;
wire [3:0] vns_videooverlaysoc_shared_sel;
wire vns_videooverlaysoc_shared_cyc;
wire vns_videooverlaysoc_shared_stb;
reg vns_videooverlaysoc_shared_ack = 1'd0;
wire vns_videooverlaysoc_shared_we;
wire [2:0] vns_videooverlaysoc_shared_cti;
wire [1:0] vns_videooverlaysoc_shared_bte;
wire vns_videooverlaysoc_shared_err;
wire [2:0] vns_videooverlaysoc_request;
reg [1:0] vns_videooverlaysoc_grant = 2'd0;
reg [4:0] vns_videooverlaysoc_slave_sel = 5'd0;
reg [4:0] vns_videooverlaysoc_slave_sel_r = 5'd0;
reg vns_videooverlaysoc_error = 1'd0;
wire vns_videooverlaysoc_wait;
wire vns_videooverlaysoc_done;
reg [16:0] vns_videooverlaysoc_count = 17'd65536;
wire [13:0] vns_videooverlaysoc_interface0_bank_bus_adr;
wire vns_videooverlaysoc_interface0_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface0_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface0_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank0_scratch3_re;
wire [7:0] vns_videooverlaysoc_csrbank0_scratch3_r;
wire [7:0] vns_videooverlaysoc_csrbank0_scratch3_w;
wire vns_videooverlaysoc_csrbank0_scratch2_re;
wire [7:0] vns_videooverlaysoc_csrbank0_scratch2_r;
wire [7:0] vns_videooverlaysoc_csrbank0_scratch2_w;
wire vns_videooverlaysoc_csrbank0_scratch1_re;
wire [7:0] vns_videooverlaysoc_csrbank0_scratch1_r;
wire [7:0] vns_videooverlaysoc_csrbank0_scratch1_w;
wire vns_videooverlaysoc_csrbank0_scratch0_re;
wire [7:0] vns_videooverlaysoc_csrbank0_scratch0_r;
wire [7:0] vns_videooverlaysoc_csrbank0_scratch0_w;
wire vns_videooverlaysoc_csrbank0_bus_errors3_re;
wire [7:0] vns_videooverlaysoc_csrbank0_bus_errors3_r;
wire [7:0] vns_videooverlaysoc_csrbank0_bus_errors3_w;
wire vns_videooverlaysoc_csrbank0_bus_errors2_re;
wire [7:0] vns_videooverlaysoc_csrbank0_bus_errors2_r;
wire [7:0] vns_videooverlaysoc_csrbank0_bus_errors2_w;
wire vns_videooverlaysoc_csrbank0_bus_errors1_re;
wire [7:0] vns_videooverlaysoc_csrbank0_bus_errors1_r;
wire [7:0] vns_videooverlaysoc_csrbank0_bus_errors1_w;
wire vns_videooverlaysoc_csrbank0_bus_errors0_re;
wire [7:0] vns_videooverlaysoc_csrbank0_bus_errors0_r;
wire [7:0] vns_videooverlaysoc_csrbank0_bus_errors0_w;
wire vns_videooverlaysoc_csrbank0_sel;
wire [13:0] vns_videooverlaysoc_interface1_bank_bus_adr;
wire vns_videooverlaysoc_interface1_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface1_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface1_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank1_half_sys8x_taps0_re;
wire [3:0] vns_videooverlaysoc_csrbank1_half_sys8x_taps0_r;
wire [3:0] vns_videooverlaysoc_csrbank1_half_sys8x_taps0_w;
wire vns_videooverlaysoc_csrbank1_dly_sel0_re;
wire [3:0] vns_videooverlaysoc_csrbank1_dly_sel0_r;
wire [3:0] vns_videooverlaysoc_csrbank1_dly_sel0_w;
wire vns_videooverlaysoc_csrbank1_sel;
wire [13:0] vns_videooverlaysoc_interface2_bank_bus_adr;
wire vns_videooverlaysoc_interface2_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface2_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface2_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank2_Km6_re;
wire [7:0] vns_videooverlaysoc_csrbank2_Km6_r;
wire [7:0] vns_videooverlaysoc_csrbank2_Km6_w;
wire vns_videooverlaysoc_csrbank2_Km5_re;
wire [7:0] vns_videooverlaysoc_csrbank2_Km5_r;
wire [7:0] vns_videooverlaysoc_csrbank2_Km5_w;
wire vns_videooverlaysoc_csrbank2_Km4_re;
wire [7:0] vns_videooverlaysoc_csrbank2_Km4_r;
wire [7:0] vns_videooverlaysoc_csrbank2_Km4_w;
wire vns_videooverlaysoc_csrbank2_Km3_re;
wire [7:0] vns_videooverlaysoc_csrbank2_Km3_r;
wire [7:0] vns_videooverlaysoc_csrbank2_Km3_w;
wire vns_videooverlaysoc_csrbank2_Km2_re;
wire [7:0] vns_videooverlaysoc_csrbank2_Km2_r;
wire [7:0] vns_videooverlaysoc_csrbank2_Km2_w;
wire vns_videooverlaysoc_csrbank2_Km1_re;
wire [7:0] vns_videooverlaysoc_csrbank2_Km1_r;
wire [7:0] vns_videooverlaysoc_csrbank2_Km1_w;
wire vns_videooverlaysoc_csrbank2_Km0_re;
wire [7:0] vns_videooverlaysoc_csrbank2_Km0_r;
wire [7:0] vns_videooverlaysoc_csrbank2_Km0_w;
wire vns_videooverlaysoc_csrbank2_Km_valid0_re;
wire vns_videooverlaysoc_csrbank2_Km_valid0_r;
wire vns_videooverlaysoc_csrbank2_Km_valid0_w;
wire vns_videooverlaysoc_csrbank2_hpd_ena0_re;
wire vns_videooverlaysoc_csrbank2_hpd_ena0_r;
wire vns_videooverlaysoc_csrbank2_hpd_ena0_w;
wire vns_videooverlaysoc_csrbank2_sel;
wire [13:0] vns_videooverlaysoc_interface3_bank_bus_adr;
wire vns_videooverlaysoc_interface3_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface3_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface3_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank3_underflow_enable0_re;
wire vns_videooverlaysoc_csrbank3_underflow_enable0_r;
wire vns_videooverlaysoc_csrbank3_underflow_enable0_w;
wire vns_videooverlaysoc_csrbank3_underflow_counter3_re;
wire [7:0] vns_videooverlaysoc_csrbank3_underflow_counter3_r;
wire [7:0] vns_videooverlaysoc_csrbank3_underflow_counter3_w;
wire vns_videooverlaysoc_csrbank3_underflow_counter2_re;
wire [7:0] vns_videooverlaysoc_csrbank3_underflow_counter2_r;
wire [7:0] vns_videooverlaysoc_csrbank3_underflow_counter2_w;
wire vns_videooverlaysoc_csrbank3_underflow_counter1_re;
wire [7:0] vns_videooverlaysoc_csrbank3_underflow_counter1_r;
wire [7:0] vns_videooverlaysoc_csrbank3_underflow_counter1_w;
wire vns_videooverlaysoc_csrbank3_underflow_counter0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_underflow_counter0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_underflow_counter0_w;
wire vns_videooverlaysoc_csrbank3_initiator_enable0_re;
wire vns_videooverlaysoc_csrbank3_initiator_enable0_r;
wire vns_videooverlaysoc_csrbank3_initiator_enable0_w;
reg [3:0] vns_videooverlaysoc_csrbank3_initiator_hres_backstore = 4'd0;
wire vns_videooverlaysoc_csrbank3_initiator_hres1_re;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_hres1_r;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_hres1_w;
wire vns_videooverlaysoc_csrbank3_initiator_hres0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_hres0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_hres0_w;
reg [3:0] vns_videooverlaysoc_csrbank3_initiator_hsync_start_backstore = 4'd0;
wire vns_videooverlaysoc_csrbank3_initiator_hsync_start1_re;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_hsync_start1_r;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_hsync_start1_w;
wire vns_videooverlaysoc_csrbank3_initiator_hsync_start0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_hsync_start0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_hsync_start0_w;
reg [3:0] vns_videooverlaysoc_csrbank3_initiator_hsync_end_backstore = 4'd0;
wire vns_videooverlaysoc_csrbank3_initiator_hsync_end1_re;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_hsync_end1_r;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_hsync_end1_w;
wire vns_videooverlaysoc_csrbank3_initiator_hsync_end0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_hsync_end0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_hsync_end0_w;
reg [3:0] vns_videooverlaysoc_csrbank3_initiator_hscan_backstore = 4'd0;
wire vns_videooverlaysoc_csrbank3_initiator_hscan1_re;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_hscan1_r;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_hscan1_w;
wire vns_videooverlaysoc_csrbank3_initiator_hscan0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_hscan0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_hscan0_w;
reg [3:0] vns_videooverlaysoc_csrbank3_initiator_vres_backstore = 4'd0;
wire vns_videooverlaysoc_csrbank3_initiator_vres1_re;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_vres1_r;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_vres1_w;
wire vns_videooverlaysoc_csrbank3_initiator_vres0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_vres0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_vres0_w;
reg [3:0] vns_videooverlaysoc_csrbank3_initiator_vsync_start_backstore = 4'd0;
wire vns_videooverlaysoc_csrbank3_initiator_vsync_start1_re;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_vsync_start1_r;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_vsync_start1_w;
wire vns_videooverlaysoc_csrbank3_initiator_vsync_start0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_vsync_start0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_vsync_start0_w;
reg [3:0] vns_videooverlaysoc_csrbank3_initiator_vsync_end_backstore = 4'd0;
wire vns_videooverlaysoc_csrbank3_initiator_vsync_end1_re;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_vsync_end1_r;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_vsync_end1_w;
wire vns_videooverlaysoc_csrbank3_initiator_vsync_end0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_vsync_end0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_vsync_end0_w;
reg [3:0] vns_videooverlaysoc_csrbank3_initiator_vscan_backstore = 4'd0;
wire vns_videooverlaysoc_csrbank3_initiator_vscan1_re;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_vscan1_r;
wire [3:0] vns_videooverlaysoc_csrbank3_initiator_vscan1_w;
wire vns_videooverlaysoc_csrbank3_initiator_vscan0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_vscan0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_vscan0_w;
reg [23:0] vns_videooverlaysoc_csrbank3_initiator_base_backstore = 24'd0;
wire vns_videooverlaysoc_csrbank3_initiator_base3_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_base3_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_base3_w;
wire vns_videooverlaysoc_csrbank3_initiator_base2_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_base2_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_base2_w;
wire vns_videooverlaysoc_csrbank3_initiator_base1_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_base1_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_base1_w;
wire vns_videooverlaysoc_csrbank3_initiator_base0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_base0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_base0_w;
reg [23:0] vns_videooverlaysoc_csrbank3_initiator_length_backstore = 24'd0;
wire vns_videooverlaysoc_csrbank3_initiator_length3_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_length3_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_length3_w;
wire vns_videooverlaysoc_csrbank3_initiator_length2_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_length2_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_length2_w;
wire vns_videooverlaysoc_csrbank3_initiator_length1_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_length1_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_length1_w;
wire vns_videooverlaysoc_csrbank3_initiator_length0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_length0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_initiator_length0_w;
wire vns_videooverlaysoc_csrbank3_dma_delay_base3_re;
wire [7:0] vns_videooverlaysoc_csrbank3_dma_delay_base3_r;
wire [7:0] vns_videooverlaysoc_csrbank3_dma_delay_base3_w;
wire vns_videooverlaysoc_csrbank3_dma_delay_base2_re;
wire [7:0] vns_videooverlaysoc_csrbank3_dma_delay_base2_r;
wire [7:0] vns_videooverlaysoc_csrbank3_dma_delay_base2_w;
wire vns_videooverlaysoc_csrbank3_dma_delay_base1_re;
wire [7:0] vns_videooverlaysoc_csrbank3_dma_delay_base1_r;
wire [7:0] vns_videooverlaysoc_csrbank3_dma_delay_base1_w;
wire vns_videooverlaysoc_csrbank3_dma_delay_base0_re;
wire [7:0] vns_videooverlaysoc_csrbank3_dma_delay_base0_r;
wire [7:0] vns_videooverlaysoc_csrbank3_dma_delay_base0_w;
wire vns_videooverlaysoc_csrbank3_sel;
wire [13:0] vns_videooverlaysoc_interface0_sram_bus_adr;
wire vns_videooverlaysoc_interface0_sram_bus_we;
wire [7:0] vns_videooverlaysoc_interface0_sram_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface0_sram_bus_dat_r = 8'd0;
wire [7:0] vns_videooverlaysoc_sram0_adr;
wire [7:0] vns_videooverlaysoc_sram0_dat_r;
wire vns_videooverlaysoc_sram0_we;
wire [7:0] vns_videooverlaysoc_sram0_dat_w;
wire vns_videooverlaysoc_sram0_sel;
reg vns_videooverlaysoc_sram0_sel_r = 1'd0;
wire [13:0] vns_videooverlaysoc_interface4_bank_bus_adr;
wire vns_videooverlaysoc_interface4_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface4_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface4_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank4_edid_hpd_notif_re;
wire vns_videooverlaysoc_csrbank4_edid_hpd_notif_r;
wire vns_videooverlaysoc_csrbank4_edid_hpd_notif_w;
wire vns_videooverlaysoc_csrbank4_edid_hpd_en0_re;
wire vns_videooverlaysoc_csrbank4_edid_hpd_en0_r;
wire vns_videooverlaysoc_csrbank4_edid_hpd_en0_w;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_reset0_re;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_reset0_r;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_reset0_w;
wire vns_videooverlaysoc_csrbank4_clocking_locked_re;
wire vns_videooverlaysoc_csrbank4_clocking_locked_r;
wire vns_videooverlaysoc_csrbank4_clocking_locked_w;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_re;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_r;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_w;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_adr0_re;
wire [6:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_adr0_r;
wire [6:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_adr0_w;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w1_re;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w1_r;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w1_w;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w0_re;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w0_r;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w0_w;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r1_re;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r1_r;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r1_w;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r0_re;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r0_r;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r0_w;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r1_re;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r1_r;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r1_w;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r0_re;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r0_r;
wire [7:0] vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r0_w;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_o_re;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_o_r;
wire vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_o_w;
wire vns_videooverlaysoc_csrbank4_data0_cap_phase_re;
wire [1:0] vns_videooverlaysoc_csrbank4_data0_cap_phase_r;
wire [1:0] vns_videooverlaysoc_csrbank4_data0_cap_phase_w;
wire vns_videooverlaysoc_csrbank4_data0_charsync_char_synced_re;
wire vns_videooverlaysoc_csrbank4_data0_charsync_char_synced_r;
wire vns_videooverlaysoc_csrbank4_data0_charsync_char_synced_w;
wire vns_videooverlaysoc_csrbank4_data0_charsync_ctl_pos_re;
wire [3:0] vns_videooverlaysoc_csrbank4_data0_charsync_ctl_pos_r;
wire [3:0] vns_videooverlaysoc_csrbank4_data0_charsync_ctl_pos_w;
wire vns_videooverlaysoc_csrbank4_data0_wer_value2_re;
wire [7:0] vns_videooverlaysoc_csrbank4_data0_wer_value2_r;
wire [7:0] vns_videooverlaysoc_csrbank4_data0_wer_value2_w;
wire vns_videooverlaysoc_csrbank4_data0_wer_value1_re;
wire [7:0] vns_videooverlaysoc_csrbank4_data0_wer_value1_r;
wire [7:0] vns_videooverlaysoc_csrbank4_data0_wer_value1_w;
wire vns_videooverlaysoc_csrbank4_data0_wer_value0_re;
wire [7:0] vns_videooverlaysoc_csrbank4_data0_wer_value0_r;
wire [7:0] vns_videooverlaysoc_csrbank4_data0_wer_value0_w;
wire vns_videooverlaysoc_csrbank4_data1_cap_phase_re;
wire [1:0] vns_videooverlaysoc_csrbank4_data1_cap_phase_r;
wire [1:0] vns_videooverlaysoc_csrbank4_data1_cap_phase_w;
wire vns_videooverlaysoc_csrbank4_data1_charsync_char_synced_re;
wire vns_videooverlaysoc_csrbank4_data1_charsync_char_synced_r;
wire vns_videooverlaysoc_csrbank4_data1_charsync_char_synced_w;
wire vns_videooverlaysoc_csrbank4_data1_charsync_ctl_pos_re;
wire [3:0] vns_videooverlaysoc_csrbank4_data1_charsync_ctl_pos_r;
wire [3:0] vns_videooverlaysoc_csrbank4_data1_charsync_ctl_pos_w;
wire vns_videooverlaysoc_csrbank4_data1_wer_value2_re;
wire [7:0] vns_videooverlaysoc_csrbank4_data1_wer_value2_r;
wire [7:0] vns_videooverlaysoc_csrbank4_data1_wer_value2_w;
wire vns_videooverlaysoc_csrbank4_data1_wer_value1_re;
wire [7:0] vns_videooverlaysoc_csrbank4_data1_wer_value1_r;
wire [7:0] vns_videooverlaysoc_csrbank4_data1_wer_value1_w;
wire vns_videooverlaysoc_csrbank4_data1_wer_value0_re;
wire [7:0] vns_videooverlaysoc_csrbank4_data1_wer_value0_r;
wire [7:0] vns_videooverlaysoc_csrbank4_data1_wer_value0_w;
wire vns_videooverlaysoc_csrbank4_data2_cap_phase_re;
wire [1:0] vns_videooverlaysoc_csrbank4_data2_cap_phase_r;
wire [1:0] vns_videooverlaysoc_csrbank4_data2_cap_phase_w;
wire vns_videooverlaysoc_csrbank4_data2_charsync_char_synced_re;
wire vns_videooverlaysoc_csrbank4_data2_charsync_char_synced_r;
wire vns_videooverlaysoc_csrbank4_data2_charsync_char_synced_w;
wire vns_videooverlaysoc_csrbank4_data2_charsync_ctl_pos_re;
wire [3:0] vns_videooverlaysoc_csrbank4_data2_charsync_ctl_pos_r;
wire [3:0] vns_videooverlaysoc_csrbank4_data2_charsync_ctl_pos_w;
wire vns_videooverlaysoc_csrbank4_data2_wer_value2_re;
wire [7:0] vns_videooverlaysoc_csrbank4_data2_wer_value2_r;
wire [7:0] vns_videooverlaysoc_csrbank4_data2_wer_value2_w;
wire vns_videooverlaysoc_csrbank4_data2_wer_value1_re;
wire [7:0] vns_videooverlaysoc_csrbank4_data2_wer_value1_r;
wire [7:0] vns_videooverlaysoc_csrbank4_data2_wer_value1_w;
wire vns_videooverlaysoc_csrbank4_data2_wer_value0_re;
wire [7:0] vns_videooverlaysoc_csrbank4_data2_wer_value0_r;
wire [7:0] vns_videooverlaysoc_csrbank4_data2_wer_value0_w;
wire vns_videooverlaysoc_csrbank4_chansync_channels_synced_re;
wire vns_videooverlaysoc_csrbank4_chansync_channels_synced_r;
wire vns_videooverlaysoc_csrbank4_chansync_channels_synced_w;
wire vns_videooverlaysoc_csrbank4_decode_terc4_dvimode0_re;
wire vns_videooverlaysoc_csrbank4_decode_terc4_dvimode0_r;
wire vns_videooverlaysoc_csrbank4_decode_terc4_dvimode0_w;
wire vns_videooverlaysoc_csrbank4_resdetection_hres1_re;
wire [2:0] vns_videooverlaysoc_csrbank4_resdetection_hres1_r;
wire [2:0] vns_videooverlaysoc_csrbank4_resdetection_hres1_w;
wire vns_videooverlaysoc_csrbank4_resdetection_hres0_re;
wire [7:0] vns_videooverlaysoc_csrbank4_resdetection_hres0_r;
wire [7:0] vns_videooverlaysoc_csrbank4_resdetection_hres0_w;
wire vns_videooverlaysoc_csrbank4_resdetection_vres1_re;
wire [2:0] vns_videooverlaysoc_csrbank4_resdetection_vres1_r;
wire [2:0] vns_videooverlaysoc_csrbank4_resdetection_vres1_w;
wire vns_videooverlaysoc_csrbank4_resdetection_vres0_re;
wire [7:0] vns_videooverlaysoc_csrbank4_resdetection_vres0_r;
wire [7:0] vns_videooverlaysoc_csrbank4_resdetection_vres0_w;
wire vns_videooverlaysoc_csrbank4_sel;
wire [13:0] vns_videooverlaysoc_interface5_bank_bus_adr;
wire vns_videooverlaysoc_interface5_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface5_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface5_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank5_value3_re;
wire [7:0] vns_videooverlaysoc_csrbank5_value3_r;
wire [7:0] vns_videooverlaysoc_csrbank5_value3_w;
wire vns_videooverlaysoc_csrbank5_value2_re;
wire [7:0] vns_videooverlaysoc_csrbank5_value2_r;
wire [7:0] vns_videooverlaysoc_csrbank5_value2_w;
wire vns_videooverlaysoc_csrbank5_value1_re;
wire [7:0] vns_videooverlaysoc_csrbank5_value1_r;
wire [7:0] vns_videooverlaysoc_csrbank5_value1_w;
wire vns_videooverlaysoc_csrbank5_value0_re;
wire [7:0] vns_videooverlaysoc_csrbank5_value0_r;
wire [7:0] vns_videooverlaysoc_csrbank5_value0_w;
wire vns_videooverlaysoc_csrbank5_sel;
wire [13:0] vns_videooverlaysoc_interface1_sram_bus_adr;
wire vns_videooverlaysoc_interface1_sram_bus_we;
wire [7:0] vns_videooverlaysoc_interface1_sram_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface1_sram_bus_dat_r = 8'd0;
wire [7:0] vns_videooverlaysoc_sram1_adr;
wire [7:0] vns_videooverlaysoc_sram1_dat_r;
wire vns_videooverlaysoc_sram1_we;
wire [7:0] vns_videooverlaysoc_sram1_dat_w;
wire vns_videooverlaysoc_sram1_sel;
reg vns_videooverlaysoc_sram1_sel_r = 1'd0;
wire [13:0] vns_videooverlaysoc_interface6_bank_bus_adr;
wire vns_videooverlaysoc_interface6_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface6_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface6_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank6_edid_hpd_notif_re;
wire vns_videooverlaysoc_csrbank6_edid_hpd_notif_r;
wire vns_videooverlaysoc_csrbank6_edid_hpd_notif_w;
wire vns_videooverlaysoc_csrbank6_edid_hpd_en0_re;
wire vns_videooverlaysoc_csrbank6_edid_hpd_en0_r;
wire vns_videooverlaysoc_csrbank6_edid_hpd_en0_w;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_reset0_re;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_reset0_r;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_reset0_w;
wire vns_videooverlaysoc_csrbank6_clocking_locked_re;
wire vns_videooverlaysoc_csrbank6_clocking_locked_r;
wire vns_videooverlaysoc_csrbank6_clocking_locked_w;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_drdy_re;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_drdy_r;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_drdy_w;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_adr0_re;
wire [6:0] vns_videooverlaysoc_csrbank6_clocking_mmcm_adr0_r;
wire [6:0] vns_videooverlaysoc_csrbank6_clocking_mmcm_adr0_w;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w1_re;
wire [7:0] vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w1_r;
wire [7:0] vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w1_w;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w0_re;
wire [7:0] vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w0_r;
wire [7:0] vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w0_w;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r1_re;
wire [7:0] vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r1_r;
wire [7:0] vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r1_w;
wire vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r0_re;
wire [7:0] vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r0_r;
wire [7:0] vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r0_w;
wire vns_videooverlaysoc_csrbank6_data0_cap_phase_re;
wire [1:0] vns_videooverlaysoc_csrbank6_data0_cap_phase_r;
wire [1:0] vns_videooverlaysoc_csrbank6_data0_cap_phase_w;
wire vns_videooverlaysoc_csrbank6_data0_charsync_char_synced_re;
wire vns_videooverlaysoc_csrbank6_data0_charsync_char_synced_r;
wire vns_videooverlaysoc_csrbank6_data0_charsync_char_synced_w;
wire vns_videooverlaysoc_csrbank6_data0_charsync_ctl_pos_re;
wire [3:0] vns_videooverlaysoc_csrbank6_data0_charsync_ctl_pos_r;
wire [3:0] vns_videooverlaysoc_csrbank6_data0_charsync_ctl_pos_w;
wire vns_videooverlaysoc_csrbank6_data0_wer_value2_re;
wire [7:0] vns_videooverlaysoc_csrbank6_data0_wer_value2_r;
wire [7:0] vns_videooverlaysoc_csrbank6_data0_wer_value2_w;
wire vns_videooverlaysoc_csrbank6_data0_wer_value1_re;
wire [7:0] vns_videooverlaysoc_csrbank6_data0_wer_value1_r;
wire [7:0] vns_videooverlaysoc_csrbank6_data0_wer_value1_w;
wire vns_videooverlaysoc_csrbank6_data0_wer_value0_re;
wire [7:0] vns_videooverlaysoc_csrbank6_data0_wer_value0_r;
wire [7:0] vns_videooverlaysoc_csrbank6_data0_wer_value0_w;
wire vns_videooverlaysoc_csrbank6_data1_cap_phase_re;
wire [1:0] vns_videooverlaysoc_csrbank6_data1_cap_phase_r;
wire [1:0] vns_videooverlaysoc_csrbank6_data1_cap_phase_w;
wire vns_videooverlaysoc_csrbank6_data1_charsync_char_synced_re;
wire vns_videooverlaysoc_csrbank6_data1_charsync_char_synced_r;
wire vns_videooverlaysoc_csrbank6_data1_charsync_char_synced_w;
wire vns_videooverlaysoc_csrbank6_data1_charsync_ctl_pos_re;
wire [3:0] vns_videooverlaysoc_csrbank6_data1_charsync_ctl_pos_r;
wire [3:0] vns_videooverlaysoc_csrbank6_data1_charsync_ctl_pos_w;
wire vns_videooverlaysoc_csrbank6_data1_wer_value2_re;
wire [7:0] vns_videooverlaysoc_csrbank6_data1_wer_value2_r;
wire [7:0] vns_videooverlaysoc_csrbank6_data1_wer_value2_w;
wire vns_videooverlaysoc_csrbank6_data1_wer_value1_re;
wire [7:0] vns_videooverlaysoc_csrbank6_data1_wer_value1_r;
wire [7:0] vns_videooverlaysoc_csrbank6_data1_wer_value1_w;
wire vns_videooverlaysoc_csrbank6_data1_wer_value0_re;
wire [7:0] vns_videooverlaysoc_csrbank6_data1_wer_value0_r;
wire [7:0] vns_videooverlaysoc_csrbank6_data1_wer_value0_w;
wire vns_videooverlaysoc_csrbank6_data2_cap_phase_re;
wire [1:0] vns_videooverlaysoc_csrbank6_data2_cap_phase_r;
wire [1:0] vns_videooverlaysoc_csrbank6_data2_cap_phase_w;
wire vns_videooverlaysoc_csrbank6_data2_charsync_char_synced_re;
wire vns_videooverlaysoc_csrbank6_data2_charsync_char_synced_r;
wire vns_videooverlaysoc_csrbank6_data2_charsync_char_synced_w;
wire vns_videooverlaysoc_csrbank6_data2_charsync_ctl_pos_re;
wire [3:0] vns_videooverlaysoc_csrbank6_data2_charsync_ctl_pos_r;
wire [3:0] vns_videooverlaysoc_csrbank6_data2_charsync_ctl_pos_w;
wire vns_videooverlaysoc_csrbank6_data2_wer_value2_re;
wire [7:0] vns_videooverlaysoc_csrbank6_data2_wer_value2_r;
wire [7:0] vns_videooverlaysoc_csrbank6_data2_wer_value2_w;
wire vns_videooverlaysoc_csrbank6_data2_wer_value1_re;
wire [7:0] vns_videooverlaysoc_csrbank6_data2_wer_value1_r;
wire [7:0] vns_videooverlaysoc_csrbank6_data2_wer_value1_w;
wire vns_videooverlaysoc_csrbank6_data2_wer_value0_re;
wire [7:0] vns_videooverlaysoc_csrbank6_data2_wer_value0_r;
wire [7:0] vns_videooverlaysoc_csrbank6_data2_wer_value0_w;
wire vns_videooverlaysoc_csrbank6_chansync_channels_synced_re;
wire vns_videooverlaysoc_csrbank6_chansync_channels_synced_r;
wire vns_videooverlaysoc_csrbank6_chansync_channels_synced_w;
wire vns_videooverlaysoc_csrbank6_decode_terc4_dvimode0_re;
wire vns_videooverlaysoc_csrbank6_decode_terc4_dvimode0_r;
wire vns_videooverlaysoc_csrbank6_decode_terc4_dvimode0_w;
wire vns_videooverlaysoc_csrbank6_resdetection_hres1_re;
wire [2:0] vns_videooverlaysoc_csrbank6_resdetection_hres1_r;
wire [2:0] vns_videooverlaysoc_csrbank6_resdetection_hres1_w;
wire vns_videooverlaysoc_csrbank6_resdetection_hres0_re;
wire [7:0] vns_videooverlaysoc_csrbank6_resdetection_hres0_r;
wire [7:0] vns_videooverlaysoc_csrbank6_resdetection_hres0_w;
wire vns_videooverlaysoc_csrbank6_resdetection_vres1_re;
wire [2:0] vns_videooverlaysoc_csrbank6_resdetection_vres1_r;
wire [2:0] vns_videooverlaysoc_csrbank6_resdetection_vres1_w;
wire vns_videooverlaysoc_csrbank6_resdetection_vres0_re;
wire [7:0] vns_videooverlaysoc_csrbank6_resdetection_vres0_r;
wire [7:0] vns_videooverlaysoc_csrbank6_resdetection_vres0_w;
wire vns_videooverlaysoc_csrbank6_dma_frame_size3_re;
wire [4:0] vns_videooverlaysoc_csrbank6_dma_frame_size3_r;
wire [4:0] vns_videooverlaysoc_csrbank6_dma_frame_size3_w;
wire vns_videooverlaysoc_csrbank6_dma_frame_size2_re;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_frame_size2_r;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_frame_size2_w;
wire vns_videooverlaysoc_csrbank6_dma_frame_size1_re;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_frame_size1_r;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_frame_size1_w;
wire vns_videooverlaysoc_csrbank6_dma_frame_size0_re;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_frame_size0_r;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_frame_size0_w;
wire vns_videooverlaysoc_csrbank6_dma_slot0_status0_re;
wire [1:0] vns_videooverlaysoc_csrbank6_dma_slot0_status0_r;
wire [1:0] vns_videooverlaysoc_csrbank6_dma_slot0_status0_w;
wire vns_videooverlaysoc_csrbank6_dma_slot0_address3_re;
wire [4:0] vns_videooverlaysoc_csrbank6_dma_slot0_address3_r;
wire [4:0] vns_videooverlaysoc_csrbank6_dma_slot0_address3_w;
wire vns_videooverlaysoc_csrbank6_dma_slot0_address2_re;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot0_address2_r;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot0_address2_w;
wire vns_videooverlaysoc_csrbank6_dma_slot0_address1_re;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot0_address1_r;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot0_address1_w;
wire vns_videooverlaysoc_csrbank6_dma_slot0_address0_re;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot0_address0_r;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot0_address0_w;
wire vns_videooverlaysoc_csrbank6_dma_slot1_status0_re;
wire [1:0] vns_videooverlaysoc_csrbank6_dma_slot1_status0_r;
wire [1:0] vns_videooverlaysoc_csrbank6_dma_slot1_status0_w;
wire vns_videooverlaysoc_csrbank6_dma_slot1_address3_re;
wire [4:0] vns_videooverlaysoc_csrbank6_dma_slot1_address3_r;
wire [4:0] vns_videooverlaysoc_csrbank6_dma_slot1_address3_w;
wire vns_videooverlaysoc_csrbank6_dma_slot1_address2_re;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot1_address2_r;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot1_address2_w;
wire vns_videooverlaysoc_csrbank6_dma_slot1_address1_re;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot1_address1_r;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot1_address1_w;
wire vns_videooverlaysoc_csrbank6_dma_slot1_address0_re;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot1_address0_r;
wire [7:0] vns_videooverlaysoc_csrbank6_dma_slot1_address0_w;
wire vns_videooverlaysoc_csrbank6_dma_ev_enable0_re;
wire [1:0] vns_videooverlaysoc_csrbank6_dma_ev_enable0_r;
wire [1:0] vns_videooverlaysoc_csrbank6_dma_ev_enable0_w;
wire vns_videooverlaysoc_csrbank6_sel;
wire [13:0] vns_videooverlaysoc_interface7_bank_bus_adr;
wire vns_videooverlaysoc_interface7_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface7_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface7_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank7_value3_re;
wire [7:0] vns_videooverlaysoc_csrbank7_value3_r;
wire [7:0] vns_videooverlaysoc_csrbank7_value3_w;
wire vns_videooverlaysoc_csrbank7_value2_re;
wire [7:0] vns_videooverlaysoc_csrbank7_value2_r;
wire [7:0] vns_videooverlaysoc_csrbank7_value2_w;
wire vns_videooverlaysoc_csrbank7_value1_re;
wire [7:0] vns_videooverlaysoc_csrbank7_value1_r;
wire [7:0] vns_videooverlaysoc_csrbank7_value1_w;
wire vns_videooverlaysoc_csrbank7_value0_re;
wire [7:0] vns_videooverlaysoc_csrbank7_value0_r;
wire [7:0] vns_videooverlaysoc_csrbank7_value0_w;
wire vns_videooverlaysoc_csrbank7_sel;
wire [13:0] vns_videooverlaysoc_interface8_bank_bus_adr;
wire vns_videooverlaysoc_interface8_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface8_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface8_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank8_edid_snoop_adr0_re;
wire [7:0] vns_videooverlaysoc_csrbank8_edid_snoop_adr0_r;
wire [7:0] vns_videooverlaysoc_csrbank8_edid_snoop_adr0_w;
wire vns_videooverlaysoc_csrbank8_edid_snoop_dat_re;
wire [7:0] vns_videooverlaysoc_csrbank8_edid_snoop_dat_r;
wire [7:0] vns_videooverlaysoc_csrbank8_edid_snoop_dat_w;
wire vns_videooverlaysoc_csrbank8_sel;
wire [13:0] vns_videooverlaysoc_interface2_sram_bus_adr;
wire vns_videooverlaysoc_interface2_sram_bus_we;
wire [7:0] vns_videooverlaysoc_interface2_sram_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface2_sram_bus_dat_r = 8'd0;
wire [4:0] vns_videooverlaysoc_sram2_adr;
wire [7:0] vns_videooverlaysoc_sram2_dat_r;
wire vns_videooverlaysoc_sram2_sel;
reg vns_videooverlaysoc_sram2_sel_r = 1'd0;
wire [13:0] vns_videooverlaysoc_interface9_bank_bus_adr;
wire vns_videooverlaysoc_interface9_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface9_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface9_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank9_hrect_start1_re;
wire [3:0] vns_videooverlaysoc_csrbank9_hrect_start1_r;
wire [3:0] vns_videooverlaysoc_csrbank9_hrect_start1_w;
wire vns_videooverlaysoc_csrbank9_hrect_start0_re;
wire [7:0] vns_videooverlaysoc_csrbank9_hrect_start0_r;
wire [7:0] vns_videooverlaysoc_csrbank9_hrect_start0_w;
wire vns_videooverlaysoc_csrbank9_hrect_end1_re;
wire [3:0] vns_videooverlaysoc_csrbank9_hrect_end1_r;
wire [3:0] vns_videooverlaysoc_csrbank9_hrect_end1_w;
wire vns_videooverlaysoc_csrbank9_hrect_end0_re;
wire [7:0] vns_videooverlaysoc_csrbank9_hrect_end0_r;
wire [7:0] vns_videooverlaysoc_csrbank9_hrect_end0_w;
wire vns_videooverlaysoc_csrbank9_vrect_start1_re;
wire [3:0] vns_videooverlaysoc_csrbank9_vrect_start1_r;
wire [3:0] vns_videooverlaysoc_csrbank9_vrect_start1_w;
wire vns_videooverlaysoc_csrbank9_vrect_start0_re;
wire [7:0] vns_videooverlaysoc_csrbank9_vrect_start0_r;
wire [7:0] vns_videooverlaysoc_csrbank9_vrect_start0_w;
wire vns_videooverlaysoc_csrbank9_vrect_end1_re;
wire [3:0] vns_videooverlaysoc_csrbank9_vrect_end1_r;
wire [3:0] vns_videooverlaysoc_csrbank9_vrect_end1_w;
wire vns_videooverlaysoc_csrbank9_vrect_end0_re;
wire [7:0] vns_videooverlaysoc_csrbank9_vrect_end0_r;
wire [7:0] vns_videooverlaysoc_csrbank9_vrect_end0_w;
wire vns_videooverlaysoc_csrbank9_rect_thresh0_re;
wire [7:0] vns_videooverlaysoc_csrbank9_rect_thresh0_r;
wire [7:0] vns_videooverlaysoc_csrbank9_rect_thresh0_w;
wire vns_videooverlaysoc_csrbank9_sel;
wire [13:0] vns_videooverlaysoc_interface10_bank_bus_adr;
wire vns_videooverlaysoc_interface10_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface10_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface10_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank10_dfii_control0_re;
wire [3:0] vns_videooverlaysoc_csrbank10_dfii_control0_r;
wire [3:0] vns_videooverlaysoc_csrbank10_dfii_control0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_command0_re;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi0_command0_r;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi0_command0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_address1_re;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi0_address1_r;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi0_address1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_address0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_address0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_address0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_baddress0_re;
wire [2:0] vns_videooverlaysoc_csrbank10_dfii_pi0_baddress0_r;
wire [2:0] vns_videooverlaysoc_csrbank10_dfii_pi0_baddress0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata7_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata7_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata7_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata6_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata6_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata6_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata5_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata5_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata5_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata4_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata4_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata4_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata3_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata3_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata3_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata2_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata2_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata2_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata1_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata1_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_rddata7_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata7_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata7_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_rddata6_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata6_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata6_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_rddata5_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata5_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata5_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_rddata4_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata4_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata4_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_rddata3_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata3_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata3_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_rddata2_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata2_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata2_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_rddata1_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata1_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi0_rddata0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi0_rddata0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_command0_re;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi1_command0_r;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi1_command0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_address1_re;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi1_address1_r;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi1_address1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_address0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_address0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_address0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_baddress0_re;
wire [2:0] vns_videooverlaysoc_csrbank10_dfii_pi1_baddress0_r;
wire [2:0] vns_videooverlaysoc_csrbank10_dfii_pi1_baddress0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata7_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata7_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata7_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata6_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata6_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata6_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata5_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata5_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata5_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata4_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata4_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata4_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata3_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata3_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata3_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata2_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata2_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata2_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata1_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata1_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_rddata7_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata7_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata7_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_rddata6_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata6_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata6_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_rddata5_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata5_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata5_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_rddata4_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata4_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata4_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_rddata3_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata3_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata3_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_rddata2_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata2_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata2_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_rddata1_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata1_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi1_rddata0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi1_rddata0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_command0_re;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi2_command0_r;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi2_command0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_address1_re;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi2_address1_r;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi2_address1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_address0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_address0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_address0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_baddress0_re;
wire [2:0] vns_videooverlaysoc_csrbank10_dfii_pi2_baddress0_r;
wire [2:0] vns_videooverlaysoc_csrbank10_dfii_pi2_baddress0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata7_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata7_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata7_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata6_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata6_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata6_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata5_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata5_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata5_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata4_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata4_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata4_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata3_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata3_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata3_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata2_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata2_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata2_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata1_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata1_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_rddata7_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata7_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata7_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_rddata6_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata6_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata6_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_rddata5_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata5_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata5_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_rddata4_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata4_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata4_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_rddata3_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata3_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata3_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_rddata2_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata2_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata2_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_rddata1_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata1_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi2_rddata0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi2_rddata0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_command0_re;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi3_command0_r;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi3_command0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_address1_re;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi3_address1_r;
wire [5:0] vns_videooverlaysoc_csrbank10_dfii_pi3_address1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_address0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_address0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_address0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_baddress0_re;
wire [2:0] vns_videooverlaysoc_csrbank10_dfii_pi3_baddress0_r;
wire [2:0] vns_videooverlaysoc_csrbank10_dfii_pi3_baddress0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata7_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata7_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata7_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata6_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata6_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata6_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata5_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata5_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata5_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata4_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata4_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata4_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata3_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata3_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata3_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata2_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata2_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata2_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata1_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata1_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata0_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_rddata7_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata7_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata7_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_rddata6_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata6_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata6_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_rddata5_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata5_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata5_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_rddata4_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata4_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata4_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_rddata3_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata3_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata3_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_rddata2_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata2_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata2_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_rddata1_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata1_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata1_w;
wire vns_videooverlaysoc_csrbank10_dfii_pi3_rddata0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_dfii_pi3_rddata0_w;
wire vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads2_re;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads2_r;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads2_w;
wire vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads1_re;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads1_r;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads1_w;
wire vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads0_w;
wire vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites2_re;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites2_r;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites2_w;
wire vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites1_re;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites1_r;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites1_w;
wire vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites0_w;
wire vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width1_re;
wire vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width1_r;
wire vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width1_w;
wire vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width0_re;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width0_r;
wire [7:0] vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width0_w;
wire vns_videooverlaysoc_csrbank10_sel;
wire [13:0] vns_videooverlaysoc_interface11_bank_bus_adr;
wire vns_videooverlaysoc_interface11_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface11_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface11_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank11_load3_re;
wire [7:0] vns_videooverlaysoc_csrbank11_load3_r;
wire [7:0] vns_videooverlaysoc_csrbank11_load3_w;
wire vns_videooverlaysoc_csrbank11_load2_re;
wire [7:0] vns_videooverlaysoc_csrbank11_load2_r;
wire [7:0] vns_videooverlaysoc_csrbank11_load2_w;
wire vns_videooverlaysoc_csrbank11_load1_re;
wire [7:0] vns_videooverlaysoc_csrbank11_load1_r;
wire [7:0] vns_videooverlaysoc_csrbank11_load1_w;
wire vns_videooverlaysoc_csrbank11_load0_re;
wire [7:0] vns_videooverlaysoc_csrbank11_load0_r;
wire [7:0] vns_videooverlaysoc_csrbank11_load0_w;
wire vns_videooverlaysoc_csrbank11_reload3_re;
wire [7:0] vns_videooverlaysoc_csrbank11_reload3_r;
wire [7:0] vns_videooverlaysoc_csrbank11_reload3_w;
wire vns_videooverlaysoc_csrbank11_reload2_re;
wire [7:0] vns_videooverlaysoc_csrbank11_reload2_r;
wire [7:0] vns_videooverlaysoc_csrbank11_reload2_w;
wire vns_videooverlaysoc_csrbank11_reload1_re;
wire [7:0] vns_videooverlaysoc_csrbank11_reload1_r;
wire [7:0] vns_videooverlaysoc_csrbank11_reload1_w;
wire vns_videooverlaysoc_csrbank11_reload0_re;
wire [7:0] vns_videooverlaysoc_csrbank11_reload0_r;
wire [7:0] vns_videooverlaysoc_csrbank11_reload0_w;
wire vns_videooverlaysoc_csrbank11_en0_re;
wire vns_videooverlaysoc_csrbank11_en0_r;
wire vns_videooverlaysoc_csrbank11_en0_w;
wire vns_videooverlaysoc_csrbank11_value3_re;
wire [7:0] vns_videooverlaysoc_csrbank11_value3_r;
wire [7:0] vns_videooverlaysoc_csrbank11_value3_w;
wire vns_videooverlaysoc_csrbank11_value2_re;
wire [7:0] vns_videooverlaysoc_csrbank11_value2_r;
wire [7:0] vns_videooverlaysoc_csrbank11_value2_w;
wire vns_videooverlaysoc_csrbank11_value1_re;
wire [7:0] vns_videooverlaysoc_csrbank11_value1_r;
wire [7:0] vns_videooverlaysoc_csrbank11_value1_w;
wire vns_videooverlaysoc_csrbank11_value0_re;
wire [7:0] vns_videooverlaysoc_csrbank11_value0_r;
wire [7:0] vns_videooverlaysoc_csrbank11_value0_w;
wire vns_videooverlaysoc_csrbank11_ev_enable0_re;
wire vns_videooverlaysoc_csrbank11_ev_enable0_r;
wire vns_videooverlaysoc_csrbank11_ev_enable0_w;
wire vns_videooverlaysoc_csrbank11_sel;
wire [13:0] vns_videooverlaysoc_interface12_bank_bus_adr;
wire vns_videooverlaysoc_interface12_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface12_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface12_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank12_txfull_re;
wire vns_videooverlaysoc_csrbank12_txfull_r;
wire vns_videooverlaysoc_csrbank12_txfull_w;
wire vns_videooverlaysoc_csrbank12_rxempty_re;
wire vns_videooverlaysoc_csrbank12_rxempty_r;
wire vns_videooverlaysoc_csrbank12_rxempty_w;
wire vns_videooverlaysoc_csrbank12_ev_enable0_re;
wire [1:0] vns_videooverlaysoc_csrbank12_ev_enable0_r;
wire [1:0] vns_videooverlaysoc_csrbank12_ev_enable0_w;
wire vns_videooverlaysoc_csrbank12_sel;
wire [13:0] vns_videooverlaysoc_interface13_bank_bus_adr;
wire vns_videooverlaysoc_interface13_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface13_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface13_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank13_tuning_word3_re;
wire [7:0] vns_videooverlaysoc_csrbank13_tuning_word3_r;
wire [7:0] vns_videooverlaysoc_csrbank13_tuning_word3_w;
wire vns_videooverlaysoc_csrbank13_tuning_word2_re;
wire [7:0] vns_videooverlaysoc_csrbank13_tuning_word2_r;
wire [7:0] vns_videooverlaysoc_csrbank13_tuning_word2_w;
wire vns_videooverlaysoc_csrbank13_tuning_word1_re;
wire [7:0] vns_videooverlaysoc_csrbank13_tuning_word1_r;
wire [7:0] vns_videooverlaysoc_csrbank13_tuning_word1_w;
wire vns_videooverlaysoc_csrbank13_tuning_word0_re;
wire [7:0] vns_videooverlaysoc_csrbank13_tuning_word0_r;
wire [7:0] vns_videooverlaysoc_csrbank13_tuning_word0_w;
wire vns_videooverlaysoc_csrbank13_sel;
wire [13:0] vns_videooverlaysoc_interface14_bank_bus_adr;
wire vns_videooverlaysoc_interface14_bank_bus_we;
wire [7:0] vns_videooverlaysoc_interface14_bank_bus_dat_w;
reg [7:0] vns_videooverlaysoc_interface14_bank_bus_dat_r = 8'd0;
wire vns_videooverlaysoc_csrbank14_temperature1_re;
wire [3:0] vns_videooverlaysoc_csrbank14_temperature1_r;
wire [3:0] vns_videooverlaysoc_csrbank14_temperature1_w;
wire vns_videooverlaysoc_csrbank14_temperature0_re;
wire [7:0] vns_videooverlaysoc_csrbank14_temperature0_r;
wire [7:0] vns_videooverlaysoc_csrbank14_temperature0_w;
wire vns_videooverlaysoc_csrbank14_vccint1_re;
wire [3:0] vns_videooverlaysoc_csrbank14_vccint1_r;
wire [3:0] vns_videooverlaysoc_csrbank14_vccint1_w;
wire vns_videooverlaysoc_csrbank14_vccint0_re;
wire [7:0] vns_videooverlaysoc_csrbank14_vccint0_r;
wire [7:0] vns_videooverlaysoc_csrbank14_vccint0_w;
wire vns_videooverlaysoc_csrbank14_vccaux1_re;
wire [3:0] vns_videooverlaysoc_csrbank14_vccaux1_r;
wire [3:0] vns_videooverlaysoc_csrbank14_vccaux1_w;
wire vns_videooverlaysoc_csrbank14_vccaux0_re;
wire [7:0] vns_videooverlaysoc_csrbank14_vccaux0_r;
wire [7:0] vns_videooverlaysoc_csrbank14_vccaux0_w;
wire vns_videooverlaysoc_csrbank14_vccbram1_re;
wire [3:0] vns_videooverlaysoc_csrbank14_vccbram1_r;
wire [3:0] vns_videooverlaysoc_csrbank14_vccbram1_w;
wire vns_videooverlaysoc_csrbank14_vccbram0_re;
wire [7:0] vns_videooverlaysoc_csrbank14_vccbram0_r;
wire [7:0] vns_videooverlaysoc_csrbank14_vccbram0_w;
wire vns_videooverlaysoc_csrbank14_sel;
wire [15:0] vns_slice_proxy0;
wire [15:0] vns_slice_proxy1;
wire [47:0] vns_slice_proxy2;
wire [47:0] vns_slice_proxy3;
wire [47:0] vns_slice_proxy4;
wire [47:0] vns_slice_proxy5;
wire [47:0] vns_slice_proxy6;
wire [47:0] vns_slice_proxy7;
wire [47:0] vns_slice_proxy8;
wire [47:0] vns_slice_proxy9;
wire [47:0] vns_slice_proxy10;
wire [47:0] vns_slice_proxy11;
wire [47:0] vns_slice_proxy12;
wire [47:0] vns_slice_proxy13;
wire [7:0] vns_slice_proxy14;
wire [15:0] vns_slice_proxy15;
wire [15:0] vns_slice_proxy16;
wire [15:0] vns_slice_proxy17;
wire [15:0] vns_slice_proxy18;
wire [15:0] vns_slice_proxy19;
wire [15:0] vns_slice_proxy20;
wire [7:0] vns_slice_proxy21;
wire [31:0] vns_slice_proxy22;
wire [31:0] vns_slice_proxy23;
wire [31:0] vns_slice_proxy24;
wire [31:0] vns_slice_proxy25;
wire [47:0] vns_slice_proxy26;
wire [47:0] vns_slice_proxy27;
wire [47:0] vns_slice_proxy28;
wire [47:0] vns_slice_proxy29;
wire [47:0] vns_slice_proxy30;
wire [47:0] vns_slice_proxy31;
wire [31:0] vns_slice_proxy32;
wire [31:0] vns_slice_proxy33;
wire [31:0] vns_slice_proxy34;
wire [31:0] vns_slice_proxy35;
wire [47:0] vns_slice_proxy36;
wire [47:0] vns_slice_proxy37;
wire [47:0] vns_slice_proxy38;
wire [47:0] vns_slice_proxy39;
wire [47:0] vns_slice_proxy40;
wire [47:0] vns_slice_proxy41;
wire [15:0] vns_slice_proxy42;
wire [15:0] vns_slice_proxy43;
wire [15:0] vns_slice_proxy44;
wire [15:0] vns_slice_proxy45;
wire [3:0] vns_slice_proxy46;
wire [7:0] vns_slice_proxy47;
wire [31:0] vns_slice_proxy48;
wire [31:0] vns_slice_proxy49;
wire [31:0] vns_slice_proxy50;
wire [31:0] vns_slice_proxy51;
wire [31:0] vns_slice_proxy52;
wire [31:0] vns_slice_proxy53;
wire [31:0] vns_slice_proxy54;
wire [31:0] vns_slice_proxy55;
wire [15:0] vns_slice_proxy56;
wire [15:0] vns_slice_proxy57;
wire [7:0] vns_slice_proxy58;
wire [3:0] vns_slice_proxy59;
wire [15:0] vns_slice_proxy60;
wire [15:0] vns_slice_proxy61;
wire [7:0] vns_slice_proxy62;
wire [7:0] vns_slice_proxy63;
wire [31:0] vns_slice_proxy64;
wire [31:0] vns_slice_proxy65;
wire [31:0] vns_slice_proxy66;
wire [31:0] vns_slice_proxy67;
wire [15:0] vns_slice_proxy68;
wire [15:0] vns_slice_proxy69;
wire [15:0] vns_slice_proxy70;
wire [15:0] vns_slice_proxy71;
wire [15:0] vns_slice_proxy72;
wire [15:0] vns_slice_proxy73;
wire [15:0] vns_slice_proxy74;
wire [15:0] vns_slice_proxy75;
wire [3:0] vns_slice_proxy76;
wire [15:0] vns_slice_proxy77;
wire [15:0] vns_slice_proxy78;
wire vns_slice_proxy79;
wire vns_slice_proxy80;
wire [3:0] vns_slice_proxy81;
wire vns_slice_proxy82;
wire [3:0] vns_slice_proxy83;
wire vns_slice_proxy84;
wire [7:0] vns_slice_proxy85;
wire vns_slice_proxy86;
wire vns_slice_proxy87;
wire [7:0] vns_slice_proxy88;
wire vns_slice_proxy89;
wire vns_slice_proxy90;
wire [7:0] vns_slice_proxy91;
wire vns_slice_proxy92;
reg vns_comb_rhs_array_muxed0 = 1'd0;
reg [13:0] vns_comb_rhs_array_muxed1 = 14'd0;
reg [2:0] vns_comb_rhs_array_muxed2 = 3'd0;
reg vns_comb_rhs_array_muxed3 = 1'd0;
reg vns_comb_rhs_array_muxed4 = 1'd0;
reg vns_comb_rhs_array_muxed5 = 1'd0;
reg vns_comb_t_array_muxed0 = 1'd0;
reg vns_comb_t_array_muxed1 = 1'd0;
reg vns_comb_t_array_muxed2 = 1'd0;
reg vns_comb_rhs_array_muxed6 = 1'd0;
reg [13:0] vns_comb_rhs_array_muxed7 = 14'd0;
reg [2:0] vns_comb_rhs_array_muxed8 = 3'd0;
reg vns_comb_rhs_array_muxed9 = 1'd0;
reg vns_comb_rhs_array_muxed10 = 1'd0;
reg vns_comb_rhs_array_muxed11 = 1'd0;
reg vns_comb_t_array_muxed3 = 1'd0;
reg vns_comb_t_array_muxed4 = 1'd0;
reg vns_comb_t_array_muxed5 = 1'd0;
reg [20:0] vns_comb_rhs_array_muxed12 = 21'd0;
reg vns_comb_rhs_array_muxed13 = 1'd0;
reg vns_comb_rhs_array_muxed14 = 1'd0;
reg [20:0] vns_comb_rhs_array_muxed15 = 21'd0;
reg vns_comb_rhs_array_muxed16 = 1'd0;
reg vns_comb_rhs_array_muxed17 = 1'd0;
reg [20:0] vns_comb_rhs_array_muxed18 = 21'd0;
reg vns_comb_rhs_array_muxed19 = 1'd0;
reg vns_comb_rhs_array_muxed20 = 1'd0;
reg [20:0] vns_comb_rhs_array_muxed21 = 21'd0;
reg vns_comb_rhs_array_muxed22 = 1'd0;
reg vns_comb_rhs_array_muxed23 = 1'd0;
reg [20:0] vns_comb_rhs_array_muxed24 = 21'd0;
reg vns_comb_rhs_array_muxed25 = 1'd0;
reg vns_comb_rhs_array_muxed26 = 1'd0;
reg [20:0] vns_comb_rhs_array_muxed27 = 21'd0;
reg vns_comb_rhs_array_muxed28 = 1'd0;
reg vns_comb_rhs_array_muxed29 = 1'd0;
reg [20:0] vns_comb_rhs_array_muxed30 = 21'd0;
reg vns_comb_rhs_array_muxed31 = 1'd0;
reg vns_comb_rhs_array_muxed32 = 1'd0;
reg [20:0] vns_comb_rhs_array_muxed33 = 21'd0;
reg vns_comb_rhs_array_muxed34 = 1'd0;
reg vns_comb_rhs_array_muxed35 = 1'd0;
reg [23:0] vns_comb_rhs_array_muxed36 = 24'd0;
reg vns_comb_rhs_array_muxed37 = 1'd0;
reg [29:0] vns_comb_rhs_array_muxed38 = 30'd0;
reg [31:0] vns_comb_rhs_array_muxed39 = 32'd0;
reg [3:0] vns_comb_rhs_array_muxed40 = 4'd0;
reg vns_comb_rhs_array_muxed41 = 1'd0;
reg vns_comb_rhs_array_muxed42 = 1'd0;
reg vns_comb_rhs_array_muxed43 = 1'd0;
reg [2:0] vns_comb_rhs_array_muxed44 = 3'd0;
reg [1:0] vns_comb_rhs_array_muxed45 = 2'd0;
reg [29:0] vns_comb_rhs_array_muxed46 = 30'd0;
reg [31:0] vns_comb_rhs_array_muxed47 = 32'd0;
reg [3:0] vns_comb_rhs_array_muxed48 = 4'd0;
reg vns_comb_rhs_array_muxed49 = 1'd0;
reg vns_comb_rhs_array_muxed50 = 1'd0;
reg vns_comb_rhs_array_muxed51 = 1'd0;
reg [2:0] vns_comb_rhs_array_muxed52 = 3'd0;
reg [1:0] vns_comb_rhs_array_muxed53 = 2'd0;
reg [9:0] vns_sync_f_array_muxed0 = 10'd0;
reg [9:0] vns_sync_f_array_muxed1 = 10'd0;
reg [9:0] vns_sync_f_array_muxed2 = 10'd0;
reg [2:0] vns_sync_rhs_array_muxed0 = 3'd0;
reg [13:0] vns_sync_rhs_array_muxed1 = 14'd0;
reg vns_sync_rhs_array_muxed2 = 1'd0;
reg vns_sync_rhs_array_muxed3 = 1'd0;
reg vns_sync_rhs_array_muxed4 = 1'd0;
reg vns_sync_rhs_array_muxed5 = 1'd0;
reg vns_sync_rhs_array_muxed6 = 1'd0;
reg [2:0] vns_sync_rhs_array_muxed7 = 3'd0;
reg [13:0] vns_sync_rhs_array_muxed8 = 14'd0;
reg vns_sync_rhs_array_muxed9 = 1'd0;
reg vns_sync_rhs_array_muxed10 = 1'd0;
reg vns_sync_rhs_array_muxed11 = 1'd0;
reg vns_sync_rhs_array_muxed12 = 1'd0;
reg vns_sync_rhs_array_muxed13 = 1'd0;
reg [2:0] vns_sync_rhs_array_muxed14 = 3'd0;
reg [13:0] vns_sync_rhs_array_muxed15 = 14'd0;
reg vns_sync_rhs_array_muxed16 = 1'd0;
reg vns_sync_rhs_array_muxed17 = 1'd0;
reg vns_sync_rhs_array_muxed18 = 1'd0;
reg vns_sync_rhs_array_muxed19 = 1'd0;
reg vns_sync_rhs_array_muxed20 = 1'd0;
reg [2:0] vns_sync_rhs_array_muxed21 = 3'd0;
reg [13:0] vns_sync_rhs_array_muxed22 = 14'd0;
reg vns_sync_rhs_array_muxed23 = 1'd0;
reg vns_sync_rhs_array_muxed24 = 1'd0;
reg vns_sync_rhs_array_muxed25 = 1'd0;
reg vns_sync_rhs_array_muxed26 = 1'd0;
reg vns_sync_rhs_array_muxed27 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl0_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl0_regs1 = 1'd0;
wire vns_xilinxasyncresetsynchronizerimpl0;
wire vns_xilinxasyncresetsynchronizerimpl0_rst_meta;
wire vns_xilinxasyncresetsynchronizerimpl1;
wire vns_xilinxasyncresetsynchronizerimpl1_rst_meta;
wire vns_xilinxasyncresetsynchronizerimpl2;
wire vns_xilinxasyncresetsynchronizerimpl2_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [5:0] vns_xilinxmultiregimpl1_regs0 = 6'd0;
(* async_reg = "true", dont_touch = "true" *) reg [5:0] vns_xilinxmultiregimpl1_regs1 = 6'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl2_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl2_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl3_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl3_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl4_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl4_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl5_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl5_regs1 = 1'd0;
wire vns_xilinxasyncresetsynchronizerimpl3;
wire vns_xilinxasyncresetsynchronizerimpl3_rst_meta;
wire vns_xilinxasyncresetsynchronizerimpl4;
wire vns_xilinxasyncresetsynchronizerimpl4_rst_meta;
wire vns_xilinxasyncresetsynchronizerimpl5;
wire vns_xilinxasyncresetsynchronizerimpl5_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl6_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl6_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl7_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl7_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl8_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl8_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl9_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl9_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl10_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl10_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl11_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl11_regs1 = 2'd0;
wire vns_xilinxmultiregimpl11;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl12_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl12_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl13_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl13_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl14_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl14_regs1 = 4'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl15_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl15_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl16_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl16_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl17_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl17_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl18_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl18_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl19_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl19_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl20_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl20_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl21_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl21_regs1 = 2'd0;
wire vns_xilinxmultiregimpl21;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl22_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl22_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl23_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl23_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl24_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl24_regs1 = 4'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl25_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl25_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl26_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl26_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl27_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl27_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl28_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl28_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl29_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl29_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl30_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl30_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl31_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl31_regs1 = 2'd0;
wire vns_xilinxmultiregimpl31;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl32_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl32_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl33_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl33_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl34_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl34_regs1 = 4'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl35_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl35_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl36_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl36_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl37_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl37_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl38_regs0 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl38_regs1 = 11'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl39_regs0 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl39_regs1 = 11'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [5:0] vns_xilinxmultiregimpl40_regs0 = 6'd0;
(* async_reg = "true", dont_touch = "true" *) reg [5:0] vns_xilinxmultiregimpl40_regs1 = 6'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl41_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl41_regs1 = 1'd0;
wire vns_xilinxmultiregimpl41;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl42_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl42_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl43_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl43_regs1 = 1'd0;
wire vns_xilinxasyncresetsynchronizerimpl6;
wire vns_xilinxasyncresetsynchronizerimpl6_rst_meta;
wire vns_xilinxasyncresetsynchronizerimpl7;
wire vns_xilinxasyncresetsynchronizerimpl7_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl44_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl44_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl45_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl45_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl46_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl46_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl47_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl47_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl48_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl48_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl49_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl49_regs1 = 2'd0;
wire vns_xilinxmultiregimpl49;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl50_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl50_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl51_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl51_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl52_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl52_regs1 = 4'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl53_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl53_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl54_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl54_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl55_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl55_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl56_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl56_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl57_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl57_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl58_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl58_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl59_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl59_regs1 = 2'd0;
wire vns_xilinxmultiregimpl59;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl60_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl60_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl61_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl61_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl62_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl62_regs1 = 4'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl63_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl63_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl64_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl64_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl65_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl65_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl66_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl66_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl67_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl67_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl68_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl68_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl69_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl69_regs1 = 2'd0;
wire vns_xilinxmultiregimpl69;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl70_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl70_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl71_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl71_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl72_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl72_regs1 = 4'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl73_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl73_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl74_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl74_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl75_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl75_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl76_regs0 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl76_regs1 = 11'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl77_regs0 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl77_regs1 = 11'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl78_regs0 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl78_regs1 = 11'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl79_regs0 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl79_regs1 = 11'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl80_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl80_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl81_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl81_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl82_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl82_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl83_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl83_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl84_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl84_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [4:0] vns_xilinxmultiregimpl85_regs0 = 5'd0;
(* async_reg = "true", dont_touch = "true" *) reg [4:0] vns_xilinxmultiregimpl85_regs1 = 5'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [4:0] vns_xilinxmultiregimpl86_regs0 = 5'd0;
(* async_reg = "true", dont_touch = "true" *) reg [4:0] vns_xilinxmultiregimpl86_regs1 = 5'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl87_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl87_regs1 = 2'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl88_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl88_regs1 = 2'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl89_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl89_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl90_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl90_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl91_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl91_regs1 = 1'd0;
wire vns_xilinxasyncresetsynchronizerimpl8_rst_meta;
wire vns_xilinxasyncresetsynchronizerimpl9_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl92_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl92_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl93_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl93_regs1 = 2'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl94_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl94_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl95_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl95_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl96_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl96_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl97_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl97_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl98_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl98_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl99_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl99_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl100_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl100_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl101_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl101_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl102_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl102_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl103_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl103_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl104_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl104_regs1 = 3'd0;

assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_reset = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_reset;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_reset = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_reset;
assign fpga_led00 = (soc_videooverlaysoc_videooverlaysoc_sys_led ^ soc_videooverlaysoc_videooverlaysoc_pcie_led);
assign fpga_led10 = 1'd0;
assign soc_videooverlaysoc_videooverlaysoc_sys_led = soc_videooverlaysoc_videooverlaysoc_sys_counter[26];
assign soc_videooverlaysoc_hdmi_in0_freq_clk0 = hdmi_in0_pix_clk;
assign soc_videooverlaysoc_hdmi_out0_clk_gen_data0 = soc_videooverlaysoc;
assign hdmi_sda_over_up = 1'd0;
assign hdmi_sda_over_dn = 1'd0;
assign soc_videooverlaysoc_early_line_end = (soc_videooverlaysoc_hdmi_in0_timing_payload_de & (~soc_videooverlaysoc_hdmi_in0_syncpol_de));
assign soc_videooverlaysoc_hdmi_in1_freq_clk0 = hdmi_in1_pix_clk;
assign soc_videooverlaysoc_hdmi_core_out0_source_source_ready = 1'd1;
assign soc_videooverlaysoc_hdmi_out0_rgb_payload_b = soc_videooverlaysoc_core_source_data_d[7:0];
assign soc_videooverlaysoc_hdmi_out0_rgb_payload_g = soc_videooverlaysoc_core_source_data_d[15:8];
assign soc_videooverlaysoc_hdmi_out0_rgb_payload_r = soc_videooverlaysoc_core_source_data_d[23:16];
assign soc_videooverlaysoc_hdmi_out0_rgb_valid = soc_videooverlaysoc_core_source_valid_d;
assign soc_videooverlaysoc_timing_rgb_delay_sink_valid = soc_videooverlaysoc_hdmi_out0_rgb_valid;
assign soc_videooverlaysoc_timing_rgb_delay_sink_ready = soc_videooverlaysoc_hdmi_out0_rgb_ready;
assign soc_videooverlaysoc_timing_rgb_delay_sink_first = soc_videooverlaysoc_hdmi_out0_rgb_first;
assign soc_videooverlaysoc_timing_rgb_delay_sink_last = soc_videooverlaysoc_hdmi_out0_rgb_last;
assign soc_videooverlaysoc_timing_rgb_delay_sink_payload_r = soc_videooverlaysoc_hdmi_out0_rgb_payload_r;
assign soc_videooverlaysoc_timing_rgb_delay_sink_payload_g = soc_videooverlaysoc_hdmi_out0_rgb_payload_g;
assign soc_videooverlaysoc_timing_rgb_delay_sink_payload_b = soc_videooverlaysoc_hdmi_out0_rgb_payload_b;
assign soc_videooverlaysoc_hdmi_out0_rgb_d_valid = soc_videooverlaysoc_timing_rgb_delay_source_valid;
assign soc_videooverlaysoc_hdmi_out0_rgb_d_ready = soc_videooverlaysoc_timing_rgb_delay_source_ready;
assign soc_videooverlaysoc_hdmi_out0_rgb_d_first = soc_videooverlaysoc_timing_rgb_delay_source_first;
assign soc_videooverlaysoc_hdmi_out0_rgb_d_last = soc_videooverlaysoc_timing_rgb_delay_source_last;
assign soc_videooverlaysoc_hdmi_out0_rgb_d_payload_r = soc_videooverlaysoc_timing_rgb_delay_source_payload_r;
assign soc_videooverlaysoc_hdmi_out0_rgb_d_payload_g = soc_videooverlaysoc_timing_rgb_delay_source_payload_g;
assign soc_videooverlaysoc_hdmi_out0_rgb_d_payload_b = soc_videooverlaysoc_timing_rgb_delay_source_payload_b;
assign soc_videooverlaysoc_hdcp_line_end = soc_videooverlaysoc_early_line_end;
assign hpd_en = soc_videooverlaysoc_hdcp_hpd_ena_storage;
always @(*) begin
	soc_videooverlaysoc_encoder0_d0 <= 8'd0;
	soc_videooverlaysoc_encoder1_d0 <= 8'd0;
	soc_videooverlaysoc_encoder2_d0 <= 8'd0;
	if (soc_videooverlaysoc_hdcp_Km_valid_storage) begin
		soc_videooverlaysoc_encoder0_d0 <= (soc_videooverlaysoc_hdmi_out0_rgb_payload_r ^ soc_videooverlaysoc_hdcp_cipher_stream[23:16]);
		soc_videooverlaysoc_encoder1_d0 <= (soc_videooverlaysoc_hdmi_out0_rgb_payload_g ^ soc_videooverlaysoc_hdcp_cipher_stream[15:8]);
		soc_videooverlaysoc_encoder2_d0 <= (soc_videooverlaysoc_hdmi_out0_rgb_payload_b ^ soc_videooverlaysoc_hdcp_cipher_stream[7:0]);
	end else begin
		soc_videooverlaysoc_encoder0_d0 <= soc_videooverlaysoc_hdmi_out0_rgb_payload_r;
		soc_videooverlaysoc_encoder1_d0 <= soc_videooverlaysoc_hdmi_out0_rgb_payload_g;
		soc_videooverlaysoc_encoder2_d0 <= soc_videooverlaysoc_hdmi_out0_rgb_payload_b;
	end
end
assign soc_videooverlaysoc_encoder0_de = 1'd1;
assign soc_videooverlaysoc_encoder0_c = 1'd0;
assign soc_videooverlaysoc_encoder1_de = 1'd1;
assign soc_videooverlaysoc_encoder1_c = 1'd0;
assign soc_videooverlaysoc_encoder2_de = 1'd1;
assign soc_videooverlaysoc_encoder2_c = 1'd0;
assign soc_videooverlaysoc_c0 = soc_videooverlaysoc_hdmi_in0_syncpol_c0;
assign soc_videooverlaysoc_c1 = soc_videooverlaysoc_hdmi_in0_syncpol_c1;
assign soc_videooverlaysoc_c2 = soc_videooverlaysoc_hdmi_in0_syncpol_c2;
assign soc_videooverlaysoc_rect_on0 = soc_videooverlaysoc_rect_on1;
assign soc_videooverlaysoc_rect_thresh = soc_videooverlaysoc_rect_thresh_storage;
assign fpga_led20 = soc_videooverlaysoc_hdmi_in0_locked;
assign fpga_led30 = 1'd0;
assign fpga_led50 = soc_videooverlaysoc_hdmi_in1_locked;
assign etherbone_clk = sys_clk;
assign etherbone_rst = sys_rst;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_error = vns_videooverlaysoc_error;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_interrupt <= 32'd0;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_interrupt[1] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_irq;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_interrupt[2] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_irq;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_interrupt[3] <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_irq;
end
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_reset = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_reset_reset_re;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors_status = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_adr[12:0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_dat_r = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_dat_r;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_we <= 4'd0;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_we[0] <= (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_cyc & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_stb) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_we) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_sel[0]);
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_we[1] <= (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_cyc & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_stb) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_we) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_sel[1]);
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_we[2] <= (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_cyc & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_stb) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_we) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_sel[2]);
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_we[3] <= (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_cyc & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_stb) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_we) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_sel[3]);
end
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_adr[11:0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_dat_r = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_dat_w;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_valid = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxtx_re;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_payload_data = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxtx_r;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_txfull_status = (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_ready);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_valid = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_valid;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_ready = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_first = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_first;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_last = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_last;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_payload_data = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_payload_data;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_trigger = (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_ready);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_valid = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_valid;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_ready = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_first = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_first;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_last = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_last;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_payload_data = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_payload_data;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxempty_status = (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_valid);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxtx_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_payload_data;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_ready = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_clear;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_trigger = (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_valid);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_clear <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_re & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_r[0])) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_clear <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_status_w <= 2'd0;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_status_w[0] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_status;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_status_w[1] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_status;
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_clear <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_re & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_r[1])) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_clear <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_w <= 2'd0;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_w[0] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_pending;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_w[1] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_pending;
end
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_irq = ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_w[0] & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_storage[0]) | (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_w[1] & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_storage[1]));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_status = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_trigger;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_status = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_trigger;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_din = {soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_in_last, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_in_first, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_in_payload_data};
assign {soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_out_last, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_out_first, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_out_payload_data} = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_dout;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_ready = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_writable;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_valid;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_in_first = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_first;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_in_last = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_last;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_in_payload_data = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_sink_payload_data;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_valid = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_readable;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_first = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_out_first;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_last = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_out_last;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_payload_data = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_fifo_out_payload_data;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_re = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_source_ready;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_re = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_readable & ((~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_readable) | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_re));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level1 = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level0 + soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_readable);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_adr <= 4'd0;
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_replace) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_adr <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_adr <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_produce;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_din;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_we = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_we & (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_writable | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_replace));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_do_read = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_readable & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_re);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_rdport_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_consume;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_dout = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_rdport_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_rdport_re = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_do_read;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_writable = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level0 != 5'd16);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_readable = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level0 != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_din = {soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_in_last, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_in_first, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_in_payload_data};
assign {soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_out_last, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_out_first, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_out_payload_data} = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_dout;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_ready = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_writable;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_valid;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_in_first = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_first;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_in_last = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_last;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_in_payload_data = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_sink_payload_data;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_valid = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_readable;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_first = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_out_first;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_last = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_out_last;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_payload_data = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_fifo_out_payload_data;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_re = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_source_ready;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_re = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_readable & ((~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_readable) | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_re));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level1 = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level0 + soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_readable);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_adr <= 4'd0;
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_replace) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_adr <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_adr <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_produce;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_din;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_we = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_we & (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_writable | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_replace));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_do_read = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_readable & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_re);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_rdport_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_consume;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_dout = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_rdport_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_rdport_re = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_do_read;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_writable = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level0 != 5'd16);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_readable = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level0 != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_trigger = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_status_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_status;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_clear <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_pending_re & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_pending_r)) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_clear <= 1'd1;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_pending_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_pending;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_irq = (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_pending_w & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_storage);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_status = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_trigger;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern <= 8'd85;
	if ((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_preamble | soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_postamble)) begin
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern <= 1'd0;
	end else begin
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern <= 7'd85;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data0;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data1;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data2;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data3;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data4;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data5;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data6;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data7;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data8;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data9;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data10;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data11;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data12;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data13;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data14;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data15;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data16;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data17;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data18;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data19;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data20;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data21;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data22;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data23;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data24;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data25;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data26;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data27;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data28;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data29;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data30;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_i = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data31;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[0] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[32] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[1] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[33] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[2] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[34] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[3] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[35] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[4] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[36] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[5] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[37] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[6] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[38] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[7] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[39] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[8] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[40] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[9] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[41] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[10] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[42] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[11] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[43] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[12] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[44] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[13] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[45] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[14] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[46] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[15] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[47] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[16] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[48] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[17] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[49] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[18] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[50] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[19] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[51] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[20] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[52] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[21] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[53] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[22] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[54] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[23] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[55] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[24] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[56] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[25] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[57] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[26] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[58] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[27] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[59] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[28] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[60] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[29] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[61] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[30] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[62] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o[1];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[31] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o[0];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata[63] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o[1];
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[0] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[32] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[1] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[33] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[2] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[34] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[3] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[35] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[4] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[36] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[5] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[37] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[6] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[38] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[7] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[39] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[8] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[40] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[9] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[41] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[10] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[42] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[11] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[43] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[12] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[44] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[13] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[45] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[14] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[46] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[15] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[47] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[16] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[48] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[17] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[49] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[18] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[50] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[19] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[51] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[20] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[52] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[21] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[53] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[22] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[54] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[23] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[55] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[24] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[56] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[25] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[57] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[26] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[58] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[27] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[59] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[28] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[60] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[29] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[61] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[30] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[62] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o[3];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[31] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o[2];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata[63] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o[3];
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[0] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[32] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[1] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[33] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[2] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[34] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[3] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[35] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[4] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[36] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[5] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[37] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[6] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[38] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[7] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[39] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[8] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[40] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[9] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[41] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[10] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[42] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[11] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[43] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[12] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[44] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[13] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[45] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[14] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[46] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[15] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[47] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[16] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[48] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[17] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[49] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[18] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[50] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[19] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[51] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[20] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[52] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[21] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[53] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[22] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[54] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[23] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[55] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[24] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[56] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[25] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[57] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[26] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[58] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[27] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[59] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[28] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[60] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[29] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[61] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[30] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[62] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o[5];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[31] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o[4];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata[63] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o[5];
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[0] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[32] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[1] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[33] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[2] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[34] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[3] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[35] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[4] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[36] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[5] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[37] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[6] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[38] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[7] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[39] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[8] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[40] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[9] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[41] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[10] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[42] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[11] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[43] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[12] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[44] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[13] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[45] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[14] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[46] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[15] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[47] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[16] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[48] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[17] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[49] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[18] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[50] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[19] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[51] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[20] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[52] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[21] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[53] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[22] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[54] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[23] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[55] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[24] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[56] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[25] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[57] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[26] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[58] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[27] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[59] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[28] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[60] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[29] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[61] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[30] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[62] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o[7];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[31] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o[6];
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata[63] <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o[7];
end
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe = ((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en[1] | soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en[2]) | soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en[3]);
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_preamble = (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en[1] & (~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en[2]));
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_postamble = (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en[3] & (~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en[2]));
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_address;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_bank = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_bank;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cas_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cas_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cs_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cs_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_ras_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_ras_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_we_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_we_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cke = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cke;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_odt = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_odt;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_reset_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_act_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_act_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_en = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata_en;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_mask = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata_mask;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata_en = soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata_valid = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata_valid;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_address;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_bank = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_bank;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cas_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cas_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cs_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cs_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_ras_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_ras_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_we_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_we_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cke = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cke;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_odt = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_odt;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_reset_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_act_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_act_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_en = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata_en;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_mask = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata_mask;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata_en = soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata_valid = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata_valid;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_address;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_bank = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_bank;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cas_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cas_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cs_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cs_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_ras_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_ras_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_we_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_we_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cke = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cke;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_odt = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_odt;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_reset_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_act_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_act_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_en = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata_en;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_mask = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata_mask;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata_en = soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata_valid = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata_valid;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_address;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_bank = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_bank;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cas_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cas_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cs_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cs_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_ras_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_ras_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_we_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_we_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cke = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cke;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_odt = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_odt;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_reset_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_act_n = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_act_n;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_en = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata_en;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_mask = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata_mask;
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata_en = soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata_valid = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_address = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_address;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_bank = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_bank;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_cas_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cas_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_cs_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cs_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_ras_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_ras_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_we_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_we_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_cke = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cke;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_odt = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_odt;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_reset_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_act_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_act_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_wrdata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_wrdata_en = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_wrdata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_wrdata_mask = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_wrdata_mask;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata_en = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_rddata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_rddata = soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_rddata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_address = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_address;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_bank = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_bank;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_cas_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cas_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_cs_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cs_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_ras_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_ras_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_we_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_we_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_cke = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cke;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_odt = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_odt;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_reset_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_act_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_act_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_wrdata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_wrdata_en = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_wrdata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_wrdata_mask = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_wrdata_mask;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata_en = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_rddata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_rddata = soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_rddata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_address = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_address;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_bank = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_bank;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_cas_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cas_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_cs_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cs_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_ras_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_ras_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_we_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_we_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_cke = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cke;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_odt = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_odt;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_reset_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_act_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_act_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_wrdata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_wrdata_en = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_wrdata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_wrdata_mask = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_wrdata_mask;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata_en = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_rddata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_rddata = soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_rddata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_address = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_address;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_bank = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_bank;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_cas_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cas_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_cs_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cs_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_ras_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_ras_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_we_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_we_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_cke = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cke;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_odt = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_odt;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_reset_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_act_n = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_act_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_wrdata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_wrdata_en = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_wrdata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_wrdata_mask = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_wrdata_mask;
assign soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata_en = soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_rddata_en;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_rddata = soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_rddata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata_valid;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_address <= 14'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_bank <= 3'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cas_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cs_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_ras_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_we_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cke <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_odt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_reset_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_act_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata_en <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata_mask <= 8'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata_en <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_address <= 14'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_bank <= 3'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cas_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cs_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_ras_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_we_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cke <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_odt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_reset_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_act_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata_en <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata_mask <= 8'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata_en <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_address <= 14'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_bank <= 3'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cas_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cs_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_ras_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_we_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cke <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_odt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_reset_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_act_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata_en <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata_mask <= 8'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata_en <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_address <= 14'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_bank <= 3'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cas_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cs_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_ras_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_we_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cke <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_odt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_reset_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_act_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata_en <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata_mask <= 8'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata_en <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata <= 64'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata_valid <= 1'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_storage[0]) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_address <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_address;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_bank <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_bank;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cas_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_cas_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cs_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_cs_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_ras_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_ras_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_we_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_we_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cke <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_cke;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_odt <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_odt;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_reset_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_reset_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_act_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_act_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_wrdata;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_wrdata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata_mask <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_wrdata_mask;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata;
		soc_videooverlaysoc_videooverlaysoc_sdram_slave_p0_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata_valid;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_address <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_address;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_bank <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_bank;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cas_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_cas_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cs_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_cs_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_ras_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_ras_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_we_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_we_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cke <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_cke;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_odt <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_odt;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_reset_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_reset_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_act_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_act_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_wrdata;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_wrdata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata_mask <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_wrdata_mask;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata;
		soc_videooverlaysoc_videooverlaysoc_sdram_slave_p1_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata_valid;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_address <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_address;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_bank <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_bank;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cas_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_cas_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cs_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_cs_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_ras_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_ras_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_we_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_we_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cke <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_cke;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_odt <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_odt;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_reset_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_reset_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_act_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_act_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_wrdata;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_wrdata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata_mask <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_wrdata_mask;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata;
		soc_videooverlaysoc_videooverlaysoc_sdram_slave_p2_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata_valid;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_address <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_address;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_bank <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_bank;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cas_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_cas_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cs_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_cs_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_ras_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_ras_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_we_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_we_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cke <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_cke;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_odt <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_odt;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_reset_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_reset_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_act_n <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_act_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_wrdata;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_wrdata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata_mask <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_wrdata_mask;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata;
		soc_videooverlaysoc_videooverlaysoc_sdram_slave_p3_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata_valid;
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_address <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_address;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_bank <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_bank;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cas_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cas_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cs_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cs_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_ras_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_ras_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_we_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_we_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_cke <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cke;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_odt <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_odt;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_reset_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_reset_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_act_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_act_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_wrdata;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_wrdata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_wrdata_mask <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_wrdata_mask;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p0_rddata_valid;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_address <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_address;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_bank <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_bank;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cas_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cas_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cs_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cs_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_ras_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_ras_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_we_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_we_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_cke <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cke;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_odt <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_odt;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_reset_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_reset_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_act_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_act_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_wrdata;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_wrdata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_wrdata_mask <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_wrdata_mask;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p1_rddata_valid;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_address <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_address;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_bank <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_bank;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cas_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cas_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cs_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cs_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_ras_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_ras_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_we_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_we_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_cke <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cke;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_odt <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_odt;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_reset_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_reset_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_act_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_act_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_wrdata;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_wrdata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_wrdata_mask <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_wrdata_mask;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p2_rddata_valid;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_address <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_address;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_bank <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_bank;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cas_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cas_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cs_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cs_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_ras_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_ras_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_we_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_we_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_cke <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cke;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_odt <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_odt;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_reset_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_reset_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_act_n <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_act_n;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_wrdata;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_wrdata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_wrdata_mask <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_wrdata_mask;
		soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata_en <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata_en;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_master_p3_rddata_valid;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cke = soc_videooverlaysoc_videooverlaysoc_sdram_storage[1];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cke = soc_videooverlaysoc_videooverlaysoc_sdram_storage[1];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cke = soc_videooverlaysoc_videooverlaysoc_sdram_storage[1];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cke = soc_videooverlaysoc_videooverlaysoc_sdram_storage[1];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_odt = soc_videooverlaysoc_videooverlaysoc_sdram_storage[2];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_odt = soc_videooverlaysoc_videooverlaysoc_sdram_storage[2];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_odt = soc_videooverlaysoc_videooverlaysoc_sdram_storage[2];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_odt = soc_videooverlaysoc_videooverlaysoc_sdram_storage[2];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_storage[3];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_storage[3];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_storage[3];
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_reset_n = soc_videooverlaysoc_videooverlaysoc_sdram_storage[3];
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_ras_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_we_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cas_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cs_n <= 1'd1;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_issue_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cs_n <= {1{(~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage[0])}};
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_we_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage[1]);
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cas_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage[2]);
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_ras_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage[3]);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cs_n <= {1{1'd1}};
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_we_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_cas_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_ras_n <= 1'd1;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_address = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_bank = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_wrdata_en = (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_issue_re & soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage[4]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata_en = (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_issue_re & soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage[5]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_wrdata_mask = 1'd0;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_ras_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_we_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cas_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cs_n <= 1'd1;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_issue_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cs_n <= {1{(~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage[0])}};
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_we_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage[1]);
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cas_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage[2]);
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_ras_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage[3]);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cs_n <= {1{1'd1}};
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_we_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_cas_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_ras_n <= 1'd1;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_address = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_bank = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_wrdata_en = (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_issue_re & soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage[4]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata_en = (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_issue_re & soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage[5]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_wrdata_mask = 1'd0;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_ras_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_we_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cas_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cs_n <= 1'd1;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_issue_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cs_n <= {1{(~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage[0])}};
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_we_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage[1]);
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cas_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage[2]);
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_ras_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage[3]);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cs_n <= {1{1'd1}};
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_we_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_cas_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_ras_n <= 1'd1;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_address = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_bank = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_wrdata_en = (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_issue_re & soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage[4]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata_en = (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_issue_re & soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage[5]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_wrdata_mask = 1'd0;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_ras_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_we_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cas_n <= 1'd1;
	soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cs_n <= 1'd1;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_issue_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cs_n <= {1{(~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage[0])}};
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_we_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage[1]);
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cas_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage[2]);
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_ras_n <= (~soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage[3]);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cs_n <= {1{1'd1}};
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_we_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_cas_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_ras_n <= 1'd1;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_address = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_bank = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_wrdata_en = (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_issue_re & soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage[4]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata_en = (soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_issue_re & soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage[5]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_wrdata = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage;
assign soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_wrdata_mask = 1'd0;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_valid = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_we = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_addr = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_lock;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_wdata_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_wdata_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_rdata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_rdata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_valid = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_we = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_addr = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_lock;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_wdata_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_wdata_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_rdata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_rdata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_valid = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_we = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_addr = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_lock;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_wdata_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_wdata_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_rdata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_rdata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_valid = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_we = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_addr = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_lock;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_wdata_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_wdata_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_rdata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_rdata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_valid = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_we = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_addr = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_lock;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_wdata_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_wdata_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_rdata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_rdata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_valid = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_we = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_addr = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_lock;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_wdata_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_wdata_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_rdata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_rdata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_valid = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_we = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_addr = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_lock;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_wdata_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_wdata_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_rdata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_rdata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_valid = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_we = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_addr = soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_lock;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_wdata_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_wdata_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_rdata_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_rdata_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_wait = (1'd1 & (~soc_videooverlaysoc_videooverlaysoc_sdram_done));
assign soc_videooverlaysoc_videooverlaysoc_sdram_done = (soc_videooverlaysoc_videooverlaysoc_sdram_count == 1'd0);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_seq_start <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_cmd_last <= 1'd0;
	vns_refresher_next_state <= 2'd0;
	vns_refresher_next_state <= vns_refresher_state;
	case (vns_refresher_state)
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid <= 1'd1;
			if (soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_seq_start <= 1'd1;
				vns_refresher_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_seq_done) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_cmd_last <= 1'd1;
				vns_refresher_next_state <= 1'd0;
			end else begin
				soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid <= 1'd1;
			end
		end
		default: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_done) begin
				vns_refresher_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_ready = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_wdata_ready | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_rdata_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_lock = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_valid | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_hit = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row == soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_addr[20:7]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ba = 1'd0;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_a <= 14'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_col_n_addr_sel) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_a <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_addr[20:7];
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_a <= ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_auto_precharge <<< 4'd10) | {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_write);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_open);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_open);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_auto_precharge <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_valid)) begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_addr[20:7] != soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_addr[20:7])) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_auto_precharge <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_close == 1'd0);
		end
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_din = {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_we};
assign {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_we} = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_dout;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_readable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_re = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_source_ready;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_replace) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_produce;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_dat_w = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_din;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_we = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_we & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_replace));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_do_read = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_readable & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_re);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_rdport_adr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_consume;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_dout = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_rdport_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_level != 4'd8);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_readable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_level != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_pipe_ce = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_ready | (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_valid_n));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_pipe_ce;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_valid_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_busy = (1'd0 | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_valid_n);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_first_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_last_n;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_refresh_gnt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_cas <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ras <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_we <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_open <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_read <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_close <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_write <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_wdata_ready <= 1'd0;
	vns_bankmachine0_next_state <= 4'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_rdata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_col_n_addr_sel <= 1'd0;
	vns_bankmachine0_next_state <= vns_bankmachine0_state;
	case (vns_bankmachine0_state)
		1'd1: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_ready)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready) begin
					vns_bankmachine0_next_state <= 3'd5;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ras <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_we <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_close <= 1'd1;
		end
		2'd2: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_ready)) begin
				vns_bankmachine0_next_state <= 3'd5;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_close <= 1'd1;
		end
		2'd3: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_col_n_addr_sel <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_open <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready) begin
					vns_bankmachine0_next_state <= 3'd7;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_refresh_gnt <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_close <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_refresh_req)) begin
				vns_bankmachine0_next_state <= 1'd0;
			end
		end
		3'd5: begin
			vns_bankmachine0_next_state <= 3'd6;
		end
		3'd6: begin
			vns_bankmachine0_next_state <= 2'd3;
		end
		3'd7: begin
			vns_bankmachine0_next_state <= 4'd8;
		end
		4'd8: begin
			vns_bankmachine0_next_state <= 1'd0;
		end
		default: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_refresh_req) begin
				vns_bankmachine0_next_state <= 3'd4;
			end else begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_valid) begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_opened) begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_hit) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid <= 1'd1;
							if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_we) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_wdata_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_write <= 1'd1;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_we <= 1'd1;
							end else begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_req_rdata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_read <= 1'd1;
							end
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_cas <= 1'd1;
							if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_auto_precharge)) begin
								vns_bankmachine0_next_state <= 2'd2;
							end
						end else begin
							vns_bankmachine0_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine0_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_ready = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_wdata_ready | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_rdata_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_lock = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_valid | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_hit = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row == soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_addr[20:7]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ba = 1'd1;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_a <= 14'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_col_n_addr_sel) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_a <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_addr[20:7];
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_a <= ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_auto_precharge <<< 4'd10) | {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_write);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_open);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_open);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_auto_precharge <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_valid)) begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_addr[20:7] != soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_addr[20:7])) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_auto_precharge <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_close == 1'd0);
		end
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_din = {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_we};
assign {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_we} = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_dout;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_readable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_re = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_source_ready;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_replace) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_produce;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_dat_w = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_din;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_we = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_we & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_replace));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_do_read = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_readable & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_re);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_rdport_adr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_consume;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_dout = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_rdport_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_level != 4'd8);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_readable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_level != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_pipe_ce = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_ready | (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_valid_n));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_pipe_ce;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_valid_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_busy = (1'd0 | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_valid_n);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_first_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_last_n;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_open <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_read <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_close <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_write <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_wdata_ready <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_rdata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_col_n_addr_sel <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_refresh_gnt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_cas <= 1'd0;
	vns_bankmachine1_next_state <= 4'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ras <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_we <= 1'd0;
	vns_bankmachine1_next_state <= vns_bankmachine1_state;
	case (vns_bankmachine1_state)
		1'd1: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_ready)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready) begin
					vns_bankmachine1_next_state <= 3'd5;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ras <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_we <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_close <= 1'd1;
		end
		2'd2: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_ready)) begin
				vns_bankmachine1_next_state <= 3'd5;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_close <= 1'd1;
		end
		2'd3: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_col_n_addr_sel <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_open <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready) begin
					vns_bankmachine1_next_state <= 3'd7;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_refresh_gnt <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_close <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_refresh_req)) begin
				vns_bankmachine1_next_state <= 1'd0;
			end
		end
		3'd5: begin
			vns_bankmachine1_next_state <= 3'd6;
		end
		3'd6: begin
			vns_bankmachine1_next_state <= 2'd3;
		end
		3'd7: begin
			vns_bankmachine1_next_state <= 4'd8;
		end
		4'd8: begin
			vns_bankmachine1_next_state <= 1'd0;
		end
		default: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_refresh_req) begin
				vns_bankmachine1_next_state <= 3'd4;
			end else begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_valid) begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_opened) begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_hit) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid <= 1'd1;
							if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_we) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_wdata_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_write <= 1'd1;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_we <= 1'd1;
							end else begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_req_rdata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_read <= 1'd1;
							end
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_cas <= 1'd1;
							if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_auto_precharge)) begin
								vns_bankmachine1_next_state <= 2'd2;
							end
						end else begin
							vns_bankmachine1_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine1_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_ready = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_wdata_ready | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_rdata_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_lock = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_valid | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_hit = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row == soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_addr[20:7]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ba = 2'd2;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_a <= 14'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_col_n_addr_sel) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_a <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_addr[20:7];
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_a <= ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_auto_precharge <<< 4'd10) | {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_write);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_open);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_open);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_auto_precharge <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_valid)) begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_addr[20:7] != soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_addr[20:7])) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_auto_precharge <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_close == 1'd0);
		end
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_din = {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_we};
assign {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_we} = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_dout;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_readable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_re = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_source_ready;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_replace) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_produce;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_dat_w = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_din;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_we = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_we & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_replace));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_do_read = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_readable & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_re);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_rdport_adr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_consume;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_dout = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_rdport_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_level != 4'd8);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_readable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_level != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_pipe_ce = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_ready | (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_valid_n));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_pipe_ce;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_valid_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_busy = (1'd0 | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_valid_n);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_first_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_last_n;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_cas <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ras <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_we <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_open <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_read <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_close <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_write <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_wdata_ready <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_rdata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_col_n_addr_sel <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_refresh_gnt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid <= 1'd0;
	vns_bankmachine2_next_state <= 4'd0;
	vns_bankmachine2_next_state <= vns_bankmachine2_state;
	case (vns_bankmachine2_state)
		1'd1: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_ready)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready) begin
					vns_bankmachine2_next_state <= 3'd5;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ras <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_we <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_close <= 1'd1;
		end
		2'd2: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_ready)) begin
				vns_bankmachine2_next_state <= 3'd5;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_close <= 1'd1;
		end
		2'd3: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_col_n_addr_sel <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_open <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready) begin
					vns_bankmachine2_next_state <= 3'd7;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_refresh_gnt <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_close <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_refresh_req)) begin
				vns_bankmachine2_next_state <= 1'd0;
			end
		end
		3'd5: begin
			vns_bankmachine2_next_state <= 3'd6;
		end
		3'd6: begin
			vns_bankmachine2_next_state <= 2'd3;
		end
		3'd7: begin
			vns_bankmachine2_next_state <= 4'd8;
		end
		4'd8: begin
			vns_bankmachine2_next_state <= 1'd0;
		end
		default: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_refresh_req) begin
				vns_bankmachine2_next_state <= 3'd4;
			end else begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_valid) begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_opened) begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_hit) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid <= 1'd1;
							if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_we) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_wdata_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_write <= 1'd1;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_we <= 1'd1;
							end else begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_req_rdata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_read <= 1'd1;
							end
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_cas <= 1'd1;
							if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_auto_precharge)) begin
								vns_bankmachine2_next_state <= 2'd2;
							end
						end else begin
							vns_bankmachine2_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine2_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_ready = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_wdata_ready | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_rdata_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_lock = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_valid | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_hit = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row == soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_addr[20:7]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ba = 2'd3;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_a <= 14'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_col_n_addr_sel) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_a <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_addr[20:7];
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_a <= ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_auto_precharge <<< 4'd10) | {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_write);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_open);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_open);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_auto_precharge <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_valid)) begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_addr[20:7] != soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_addr[20:7])) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_auto_precharge <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_close == 1'd0);
		end
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_din = {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_we};
assign {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_we} = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_dout;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_readable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_re = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_source_ready;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_replace) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_produce;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_dat_w = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_din;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_we = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_we & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_replace));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_do_read = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_readable & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_re);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_rdport_adr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_consume;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_dout = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_rdport_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_level != 4'd8);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_readable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_level != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_pipe_ce = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_ready | (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_valid_n));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_pipe_ce;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_valid_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_busy = (1'd0 | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_valid_n);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_first_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_last_n;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_rdata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_col_n_addr_sel <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_refresh_gnt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_close <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_cas <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ras <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_we <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_open <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_read <= 1'd0;
	vns_bankmachine3_next_state <= 4'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_write <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_wdata_ready <= 1'd0;
	vns_bankmachine3_next_state <= vns_bankmachine3_state;
	case (vns_bankmachine3_state)
		1'd1: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_ready)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready) begin
					vns_bankmachine3_next_state <= 3'd5;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ras <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_we <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_close <= 1'd1;
		end
		2'd2: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_ready)) begin
				vns_bankmachine3_next_state <= 3'd5;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_close <= 1'd1;
		end
		2'd3: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_col_n_addr_sel <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_open <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready) begin
					vns_bankmachine3_next_state <= 3'd7;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_refresh_gnt <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_close <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_refresh_req)) begin
				vns_bankmachine3_next_state <= 1'd0;
			end
		end
		3'd5: begin
			vns_bankmachine3_next_state <= 3'd6;
		end
		3'd6: begin
			vns_bankmachine3_next_state <= 2'd3;
		end
		3'd7: begin
			vns_bankmachine3_next_state <= 4'd8;
		end
		4'd8: begin
			vns_bankmachine3_next_state <= 1'd0;
		end
		default: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_refresh_req) begin
				vns_bankmachine3_next_state <= 3'd4;
			end else begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_valid) begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_opened) begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_hit) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid <= 1'd1;
							if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_we) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_wdata_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_write <= 1'd1;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_we <= 1'd1;
							end else begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_req_rdata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_read <= 1'd1;
							end
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_cas <= 1'd1;
							if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_auto_precharge)) begin
								vns_bankmachine3_next_state <= 2'd2;
							end
						end else begin
							vns_bankmachine3_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine3_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_ready = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_wdata_ready | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_rdata_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_lock = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_valid | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_hit = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row == soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_addr[20:7]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ba = 3'd4;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_a <= 14'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_col_n_addr_sel) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_a <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_addr[20:7];
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_a <= ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_auto_precharge <<< 4'd10) | {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_write);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_open);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_open);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_auto_precharge <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_valid)) begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_addr[20:7] != soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_addr[20:7])) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_auto_precharge <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_close == 1'd0);
		end
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_din = {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_we};
assign {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_we} = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_dout;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_readable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_re = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_source_ready;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_replace) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_produce;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_dat_w = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_din;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_we = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_we & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_replace));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_do_read = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_readable & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_re);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_rdport_adr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_consume;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_dout = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_rdport_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_level != 4'd8);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_readable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_level != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_pipe_ce = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_ready | (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_valid_n));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_pipe_ce;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_valid_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_busy = (1'd0 | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_valid_n);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_first_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_last_n;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ras <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_we <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_open <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_read <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_close <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_write <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_wdata_ready <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_rdata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_col_n_addr_sel <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_refresh_gnt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid <= 1'd0;
	vns_bankmachine4_next_state <= 4'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_cas <= 1'd0;
	vns_bankmachine4_next_state <= vns_bankmachine4_state;
	case (vns_bankmachine4_state)
		1'd1: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_ready)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready) begin
					vns_bankmachine4_next_state <= 3'd5;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ras <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_we <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_close <= 1'd1;
		end
		2'd2: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_ready)) begin
				vns_bankmachine4_next_state <= 3'd5;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_close <= 1'd1;
		end
		2'd3: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_col_n_addr_sel <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_open <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready) begin
					vns_bankmachine4_next_state <= 3'd7;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_refresh_gnt <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_close <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_refresh_req)) begin
				vns_bankmachine4_next_state <= 1'd0;
			end
		end
		3'd5: begin
			vns_bankmachine4_next_state <= 3'd6;
		end
		3'd6: begin
			vns_bankmachine4_next_state <= 2'd3;
		end
		3'd7: begin
			vns_bankmachine4_next_state <= 4'd8;
		end
		4'd8: begin
			vns_bankmachine4_next_state <= 1'd0;
		end
		default: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_refresh_req) begin
				vns_bankmachine4_next_state <= 3'd4;
			end else begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_valid) begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_opened) begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_hit) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid <= 1'd1;
							if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_we) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_wdata_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_write <= 1'd1;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_we <= 1'd1;
							end else begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_req_rdata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_read <= 1'd1;
							end
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_cas <= 1'd1;
							if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_auto_precharge)) begin
								vns_bankmachine4_next_state <= 2'd2;
							end
						end else begin
							vns_bankmachine4_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine4_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_ready = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_wdata_ready | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_rdata_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_lock = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_valid | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_hit = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row == soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_addr[20:7]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ba = 3'd5;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_a <= 14'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_col_n_addr_sel) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_a <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_addr[20:7];
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_a <= ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_auto_precharge <<< 4'd10) | {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_write);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_open);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_open);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_auto_precharge <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_valid)) begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_addr[20:7] != soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_addr[20:7])) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_auto_precharge <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_close == 1'd0);
		end
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_din = {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_we};
assign {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_we} = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_dout;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_readable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_re = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_source_ready;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_replace) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_produce;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_dat_w = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_din;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_we = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_we & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_replace));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_do_read = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_readable & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_re);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_rdport_adr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_consume;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_dout = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_rdport_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_level != 4'd8);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_readable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_level != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_pipe_ce = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_ready | (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_valid_n));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_pipe_ce;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_valid_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_busy = (1'd0 | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_valid_n);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_first_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_last_n;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_cas <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ras <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_we <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_open <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_read <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_close <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_write <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_wdata_ready <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_rdata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_col_n_addr_sel <= 1'd0;
	vns_bankmachine5_next_state <= 4'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_refresh_gnt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid <= 1'd0;
	vns_bankmachine5_next_state <= vns_bankmachine5_state;
	case (vns_bankmachine5_state)
		1'd1: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_ready)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready) begin
					vns_bankmachine5_next_state <= 3'd5;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ras <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_we <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_close <= 1'd1;
		end
		2'd2: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_ready)) begin
				vns_bankmachine5_next_state <= 3'd5;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_close <= 1'd1;
		end
		2'd3: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_col_n_addr_sel <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_open <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready) begin
					vns_bankmachine5_next_state <= 3'd7;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_refresh_gnt <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_close <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_refresh_req)) begin
				vns_bankmachine5_next_state <= 1'd0;
			end
		end
		3'd5: begin
			vns_bankmachine5_next_state <= 3'd6;
		end
		3'd6: begin
			vns_bankmachine5_next_state <= 2'd3;
		end
		3'd7: begin
			vns_bankmachine5_next_state <= 4'd8;
		end
		4'd8: begin
			vns_bankmachine5_next_state <= 1'd0;
		end
		default: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_refresh_req) begin
				vns_bankmachine5_next_state <= 3'd4;
			end else begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_valid) begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_opened) begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_hit) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid <= 1'd1;
							if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_we) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_wdata_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_write <= 1'd1;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_we <= 1'd1;
							end else begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_req_rdata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_read <= 1'd1;
							end
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_cas <= 1'd1;
							if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_auto_precharge)) begin
								vns_bankmachine5_next_state <= 2'd2;
							end
						end else begin
							vns_bankmachine5_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine5_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_ready = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_wdata_ready | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_rdata_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_lock = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_valid | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_hit = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row == soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_addr[20:7]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ba = 3'd6;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_a <= 14'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_col_n_addr_sel) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_a <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_addr[20:7];
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_a <= ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_auto_precharge <<< 4'd10) | {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_write);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_open);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_open);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_auto_precharge <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_valid)) begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_addr[20:7] != soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_addr[20:7])) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_auto_precharge <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_close == 1'd0);
		end
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_din = {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_we};
assign {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_we} = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_dout;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_readable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_re = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_source_ready;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_replace) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_produce;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_dat_w = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_din;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_we = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_we & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_replace));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_do_read = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_readable & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_re);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_rdport_adr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_consume;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_dout = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_rdport_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_level != 4'd8);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_readable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_level != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_pipe_ce = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_ready | (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_valid_n));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_pipe_ce;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_valid_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_busy = (1'd0 | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_valid_n);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_first_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_last_n;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_close <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_write <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_wdata_ready <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_rdata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_col_n_addr_sel <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_refresh_gnt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_cas <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ras <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_we <= 1'd0;
	vns_bankmachine6_next_state <= 4'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_open <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_read <= 1'd0;
	vns_bankmachine6_next_state <= vns_bankmachine6_state;
	case (vns_bankmachine6_state)
		1'd1: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_ready)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready) begin
					vns_bankmachine6_next_state <= 3'd5;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ras <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_we <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_close <= 1'd1;
		end
		2'd2: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_ready)) begin
				vns_bankmachine6_next_state <= 3'd5;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_close <= 1'd1;
		end
		2'd3: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_col_n_addr_sel <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_open <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready) begin
					vns_bankmachine6_next_state <= 3'd7;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_refresh_gnt <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_close <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_refresh_req)) begin
				vns_bankmachine6_next_state <= 1'd0;
			end
		end
		3'd5: begin
			vns_bankmachine6_next_state <= 3'd6;
		end
		3'd6: begin
			vns_bankmachine6_next_state <= 2'd3;
		end
		3'd7: begin
			vns_bankmachine6_next_state <= 4'd8;
		end
		4'd8: begin
			vns_bankmachine6_next_state <= 1'd0;
		end
		default: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_refresh_req) begin
				vns_bankmachine6_next_state <= 3'd4;
			end else begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_valid) begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_opened) begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_hit) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid <= 1'd1;
							if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_we) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_wdata_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_write <= 1'd1;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_we <= 1'd1;
							end else begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_req_rdata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_read <= 1'd1;
							end
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_cas <= 1'd1;
							if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_auto_precharge)) begin
								vns_bankmachine6_next_state <= 2'd2;
							end
						end else begin
							vns_bankmachine6_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine6_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_ready = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_wdata_ready | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_rdata_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_lock = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_valid | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_valid);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_hit = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row == soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_addr[20:7]);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ba = 3'd7;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_a <= 14'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_col_n_addr_sel) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_a <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_addr[20:7];
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_a <= ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_auto_precharge <<< 4'd10) | {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_write);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_open);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_open);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_auto_precharge <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_valid)) begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_addr[20:7] != soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_addr[20:7])) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_auto_precharge <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_close == 1'd0);
		end
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_din = {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_we};
assign {soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_last, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_first, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_addr, soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_we} = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_dout;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_readable;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_first;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_last;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_we = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_we;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_addr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_addr;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_re = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_source_ready;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_replace) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_produce;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_dat_w = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_din;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_we = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_we & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_replace));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_do_read = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_readable & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_re);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_rdport_adr = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_consume;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_dout = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_rdport_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_level != 4'd8);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_readable = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_level != 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_pipe_ce = (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_ready | (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_valid_n));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_ready = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_pipe_ce;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_valid = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_valid_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_busy = (1'd0 | soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_valid_n);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_first = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_first_n;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_last = soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_last_n;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_cas <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ras <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_we <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_open <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_read <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_close <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_write <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_wdata_ready <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_rdata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_col_n_addr_sel <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_refresh_gnt <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid <= 1'd0;
	vns_bankmachine7_next_state <= 4'd0;
	vns_bankmachine7_next_state <= vns_bankmachine7_state;
	case (vns_bankmachine7_state)
		1'd1: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_ready)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready) begin
					vns_bankmachine7_next_state <= 3'd5;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ras <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_we <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_close <= 1'd1;
		end
		2'd2: begin
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_ready)) begin
				vns_bankmachine7_next_state <= 3'd5;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_close <= 1'd1;
		end
		2'd3: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_col_n_addr_sel <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_open <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready) begin
					vns_bankmachine7_next_state <= 3'd7;
				end
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_ready) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_refresh_gnt <= 1'd1;
			end
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_close <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_refresh_req)) begin
				vns_bankmachine7_next_state <= 1'd0;
			end
		end
		3'd5: begin
			vns_bankmachine7_next_state <= 3'd6;
		end
		3'd6: begin
			vns_bankmachine7_next_state <= 2'd3;
		end
		3'd7: begin
			vns_bankmachine7_next_state <= 4'd8;
		end
		4'd8: begin
			vns_bankmachine7_next_state <= 1'd0;
		end
		default: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_refresh_req) begin
				vns_bankmachine7_next_state <= 3'd4;
			end else begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_valid) begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_opened) begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_hit) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid <= 1'd1;
							if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_we) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_wdata_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_write <= 1'd1;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_we <= 1'd1;
							end else begin
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_req_rdata_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready;
								soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_read <= 1'd1;
							end
							soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_cas <= 1'd1;
							if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_auto_precharge)) begin
								vns_bankmachine7_next_state <= 2'd2;
							end
						end else begin
							vns_bankmachine7_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine7_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we)));
assign soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we)));
assign soc_videooverlaysoc_videooverlaysoc_sdram_ras_allowed = (soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_ready & soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_ready);
assign soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_write | soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_read));
assign soc_videooverlaysoc_videooverlaysoc_sdram_cas_allowed = soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_ready;
assign soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_valid = ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_write);
assign soc_videooverlaysoc_videooverlaysoc_sdram_read_available = ((((((((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_read) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_read)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_read)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_read)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_read)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_read)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_read)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_read));
assign soc_videooverlaysoc_videooverlaysoc_sdram_write_available = ((((((((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_write) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_write)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_write)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_write)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_write)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_write)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_write)) | (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_write));
assign soc_videooverlaysoc_videooverlaysoc_sdram_max_time0 = (soc_videooverlaysoc_videooverlaysoc_sdram_time0 == 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_sdram_max_time1 = (soc_videooverlaysoc_videooverlaysoc_sdram_time1 == 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_refresh_req = soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_refresh_req = soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_refresh_req = soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_refresh_req = soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_refresh_req = soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_refresh_req = soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_refresh_req = soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_refresh_req = soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid;
assign soc_videooverlaysoc_videooverlaysoc_sdram_go_to_refresh = (((((((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_refresh_gnt & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_refresh_gnt) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_refresh_gnt) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_refresh_gnt) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_refresh_gnt) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_refresh_gnt) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_refresh_gnt) & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_refresh_gnt);
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_rdata = {soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_rddata, soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_rddata, soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_rddata, soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_rddata};
assign {soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_wrdata, soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_wrdata, soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_wrdata, soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_wrdata} = soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata;
assign {soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_wrdata_mask, soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_wrdata_mask, soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_wrdata_mask, soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_wrdata_mask} = (~soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata_we);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids <= 8'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[0] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[1] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[2] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[3] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[4] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[5] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[6] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[7] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_writes))));
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request = soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid = vns_comb_rhs_array_muxed0;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_a = vns_comb_rhs_array_muxed1;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ba = vns_comb_rhs_array_muxed2;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_read = vns_comb_rhs_array_muxed3;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_write = vns_comb_rhs_array_muxed4;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_cmd = vns_comb_rhs_array_muxed5;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas <= 1'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas <= vns_comb_t_array_muxed0;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras <= 1'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras <= vns_comb_t_array_muxed1;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we <= 1'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we <= vns_comb_t_array_muxed2;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_ce = (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready | (~soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid));
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids <= 8'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[0] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[1] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[2] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[3] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[4] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[5] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[6] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes))));
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[7] <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_valid & (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_cmd & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_cmds) & ((~((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_activates)) | ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_read == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads) & (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_write == soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes))));
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request = soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid = vns_comb_rhs_array_muxed6;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_a = vns_comb_rhs_array_muxed7;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ba = vns_comb_rhs_array_muxed8;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_read = vns_comb_rhs_array_muxed9;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_write = vns_comb_rhs_array_muxed10;
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_cmd = vns_comb_rhs_array_muxed11;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_cas <= 1'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_cas <= vns_comb_t_array_muxed3;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ras <= 1'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ras <= vns_comb_t_array_muxed4;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_we <= 1'd0;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_we <= vns_comb_t_array_muxed5;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant == 1'd0))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready <= 1'd1;
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant == 1'd0))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant == 1'd1))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready <= 1'd1;
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant == 1'd1))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant == 2'd2))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready <= 1'd1;
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant == 2'd2))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant == 2'd3))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready <= 1'd1;
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant == 2'd3))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant == 3'd4))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready <= 1'd1;
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant == 3'd4))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant == 3'd5))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready <= 1'd1;
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant == 3'd5))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant == 3'd6))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready <= 1'd1;
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant == 3'd6))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant == 3'd7))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready <= 1'd1;
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant == 3'd7))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_ready <= 1'd1;
	end
end
assign soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_ce = (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready | (~soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid));
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_reset_n = 1'd1;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cke = {1{soc_videooverlaysoc_videooverlaysoc_sdram_steerer0}};
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_odt = {1{soc_videooverlaysoc_videooverlaysoc_sdram_steerer1}};
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_reset_n = 1'd1;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cke = {1{soc_videooverlaysoc_videooverlaysoc_sdram_steerer2}};
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_odt = {1{soc_videooverlaysoc_videooverlaysoc_sdram_steerer3}};
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_reset_n = 1'd1;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cke = {1{soc_videooverlaysoc_videooverlaysoc_sdram_steerer4}};
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_odt = {1{soc_videooverlaysoc_videooverlaysoc_sdram_steerer5}};
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_reset_n = 1'd1;
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cke = {1{soc_videooverlaysoc_videooverlaysoc_sdram_steerer6}};
assign soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_odt = {1{soc_videooverlaysoc_videooverlaysoc_sdram_steerer7}};
assign soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_count = ((((soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_window[0] + soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_window[1]) + soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_window[2]) + soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_window[3]) + soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_window[4]);
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_en1 <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3 <= 2'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0 <= 2'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1 <= 2'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2 <= 2'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates <= 1'd0;
	vns_multiplexer_next_state <= 4'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_en0 <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready <= 1'd0;
	vns_multiplexer_next_state <= vns_multiplexer_state;
	case (vns_multiplexer_state)
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_sdram_en1 <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_writes <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates <= soc_videooverlaysoc_videooverlaysoc_sdram_ras_allowed;
			soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready <= ((~((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_ras_allowed);
			soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_cas_allowed;
			soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0 <= 1'd0;
			soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1 <= 1'd0;
			soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2 <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3 <= 2'd2;
			if (soc_videooverlaysoc_videooverlaysoc_sdram_read_available) begin
				if (((~soc_videooverlaysoc_videooverlaysoc_sdram_write_available) | soc_videooverlaysoc_videooverlaysoc_sdram_max_time1)) begin
					vns_multiplexer_next_state <= 2'd3;
				end
			end
			if (soc_videooverlaysoc_videooverlaysoc_sdram_go_to_refresh) begin
				vns_multiplexer_next_state <= 2'd2;
			end
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0 <= 2'd3;
			soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready <= 1'd1;
			if (soc_videooverlaysoc_videooverlaysoc_sdram_cmd_last) begin
				vns_multiplexer_next_state <= 1'd0;
			end
		end
		2'd3: begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_ready) begin
				vns_multiplexer_next_state <= 1'd0;
			end
		end
		3'd4: begin
			vns_multiplexer_next_state <= 3'd5;
		end
		3'd5: begin
			vns_multiplexer_next_state <= 3'd6;
		end
		3'd6: begin
			vns_multiplexer_next_state <= 3'd7;
		end
		3'd7: begin
			vns_multiplexer_next_state <= 4'd8;
		end
		4'd8: begin
			vns_multiplexer_next_state <= 4'd9;
		end
		4'd9: begin
			vns_multiplexer_next_state <= 4'd10;
		end
		4'd10: begin
			vns_multiplexer_next_state <= 4'd11;
		end
		4'd11: begin
			vns_multiplexer_next_state <= 1'd1;
		end
		default: begin
			soc_videooverlaysoc_videooverlaysoc_sdram_en0 <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_want_reads <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_want_activates <= soc_videooverlaysoc_videooverlaysoc_sdram_ras_allowed;
			soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready <= ((~((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras & (~soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas)) & (~soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we))) | soc_videooverlaysoc_videooverlaysoc_sdram_ras_allowed);
			soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_cas_allowed;
			soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0 <= 1'd0;
			soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1 <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2 <= 2'd2;
			soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3 <= 1'd0;
			if (soc_videooverlaysoc_videooverlaysoc_sdram_write_available) begin
				if (((~soc_videooverlaysoc_videooverlaysoc_sdram_read_available) | soc_videooverlaysoc_videooverlaysoc_sdram_max_time0)) begin
					vns_multiplexer_next_state <= 3'd4;
				end
			end
			if (soc_videooverlaysoc_videooverlaysoc_sdram_go_to_refresh) begin
				vns_multiplexer_next_state <= 2'd2;
			end
		end
	endcase
end
assign vns_roundrobin0_request = {(((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 1'd0) & (~(((((((vns_locked2 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid), (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 1'd0) & (~(((((((vns_locked1 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid), (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 1'd0) & (~(((((((vns_locked0 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid)};
assign vns_roundrobin0_ce = ((~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_valid) & (~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock));
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_addr = vns_comb_rhs_array_muxed12;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_we = vns_comb_rhs_array_muxed13;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_valid = vns_comb_rhs_array_muxed14;
assign vns_roundrobin1_request = {(((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 1'd1) & (~(((((((vns_locked5 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid), (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 1'd1) & (~(((((((vns_locked4 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid), (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 1'd1) & (~(((((((vns_locked3 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid)};
assign vns_roundrobin1_ce = ((~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_valid) & (~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock));
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_addr = vns_comb_rhs_array_muxed15;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_we = vns_comb_rhs_array_muxed16;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_valid = vns_comb_rhs_array_muxed17;
assign vns_roundrobin2_request = {(((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 2'd2) & (~(((((((vns_locked8 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid), (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 2'd2) & (~(((((((vns_locked7 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid), (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 2'd2) & (~(((((((vns_locked6 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid)};
assign vns_roundrobin2_ce = ((~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_valid) & (~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock));
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_addr = vns_comb_rhs_array_muxed18;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_we = vns_comb_rhs_array_muxed19;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_valid = vns_comb_rhs_array_muxed20;
assign vns_roundrobin3_request = {(((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 2'd3) & (~(((((((vns_locked11 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid), (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 2'd3) & (~(((((((vns_locked10 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid), (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 2'd3) & (~(((((((vns_locked9 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid)};
assign vns_roundrobin3_ce = ((~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_valid) & (~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock));
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_addr = vns_comb_rhs_array_muxed21;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_we = vns_comb_rhs_array_muxed22;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_valid = vns_comb_rhs_array_muxed23;
assign vns_roundrobin4_request = {(((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd4) & (~(((((((vns_locked14 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid), (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd4) & (~(((((((vns_locked13 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid), (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd4) & (~(((((((vns_locked12 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid)};
assign vns_roundrobin4_ce = ((~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_valid) & (~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock));
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_addr = vns_comb_rhs_array_muxed24;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_we = vns_comb_rhs_array_muxed25;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_valid = vns_comb_rhs_array_muxed26;
assign vns_roundrobin5_request = {(((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd5) & (~(((((((vns_locked17 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid), (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd5) & (~(((((((vns_locked16 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid), (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd5) & (~(((((((vns_locked15 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid)};
assign vns_roundrobin5_ce = ((~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_valid) & (~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock));
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_addr = vns_comb_rhs_array_muxed27;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_we = vns_comb_rhs_array_muxed28;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_valid = vns_comb_rhs_array_muxed29;
assign vns_roundrobin6_request = {(((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd6) & (~(((((((vns_locked20 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid), (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd6) & (~(((((((vns_locked19 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid), (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd6) & (~(((((((vns_locked18 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid)};
assign vns_roundrobin6_ce = ((~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_valid) & (~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock));
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_addr = vns_comb_rhs_array_muxed30;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_we = vns_comb_rhs_array_muxed31;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_valid = vns_comb_rhs_array_muxed32;
assign vns_roundrobin7_request = {(((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd7) & (~(((((((vns_locked23 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid), (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd7) & (~(((((((vns_locked22 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid), (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd7) & (~(((((((vns_locked21 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid)};
assign vns_roundrobin7_ce = ((~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_valid) & (~soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock));
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_addr = vns_comb_rhs_array_muxed33;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_we = vns_comb_rhs_array_muxed34;
assign soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_valid = vns_comb_rhs_array_muxed35;
assign soc_videooverlaysoc_videooverlaysoc_port_cmd_ready = ((((((((1'd0 | (((vns_roundrobin0_grant == 1'd0) & ((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 1'd0) & (~(((((((vns_locked0 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_ready)) | (((vns_roundrobin1_grant == 1'd0) & ((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 1'd1) & (~(((((((vns_locked3 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_ready)) | (((vns_roundrobin2_grant == 1'd0) & ((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 2'd2) & (~(((((((vns_locked6 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_ready)) | (((vns_roundrobin3_grant == 1'd0) & ((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 2'd3) & (~(((((((vns_locked9 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_ready)) | (((vns_roundrobin4_grant == 1'd0) & ((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd4) & (~(((((((vns_locked12 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_ready)) | (((vns_roundrobin5_grant == 1'd0) & ((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd5) & (~(((((((vns_locked15 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_ready)) | (((vns_roundrobin6_grant == 1'd0) & ((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd6) & (~(((((((vns_locked18 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_ready)) | (((vns_roundrobin7_grant == 1'd0) & ((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd7) & (~(((((((vns_locked21 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_ready));
assign soc_videooverlaysoc_litedramcrossbar_cmd_ready = ((((((((1'd0 | (((vns_roundrobin0_grant == 1'd1) & ((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 1'd0) & (~(((((((vns_locked1 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_ready)) | (((vns_roundrobin1_grant == 1'd1) & ((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 1'd1) & (~(((((((vns_locked4 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_ready)) | (((vns_roundrobin2_grant == 1'd1) & ((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 2'd2) & (~(((((((vns_locked7 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_ready)) | (((vns_roundrobin3_grant == 1'd1) & ((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 2'd3) & (~(((((((vns_locked10 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_ready)) | (((vns_roundrobin4_grant == 1'd1) & ((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd4) & (~(((((((vns_locked13 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_ready)) | (((vns_roundrobin5_grant == 1'd1) & ((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd5) & (~(((((((vns_locked16 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_ready)) | (((vns_roundrobin6_grant == 1'd1) & ((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd6) & (~(((((((vns_locked19 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_ready)) | (((vns_roundrobin7_grant == 1'd1) & ((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd7) & (~(((((((vns_locked22 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_ready));
assign soc_videooverlaysoc_out_dram_port_cmd_ready = ((((((((1'd0 | (((vns_roundrobin0_grant == 2'd2) & ((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 1'd0) & (~(((((((vns_locked2 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_ready)) | (((vns_roundrobin1_grant == 2'd2) & ((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 1'd1) & (~(((((((vns_locked5 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_ready)) | (((vns_roundrobin2_grant == 2'd2) & ((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 2'd2) & (~(((((((vns_locked8 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_ready)) | (((vns_roundrobin3_grant == 2'd2) & ((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 2'd3) & (~(((((((vns_locked11 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_ready)) | (((vns_roundrobin4_grant == 2'd2) & ((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd4) & (~(((((((vns_locked14 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_ready)) | (((vns_roundrobin5_grant == 2'd2) & ((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd5) & (~(((((((vns_locked17 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_ready)) | (((vns_roundrobin6_grant == 2'd2) & ((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd6) & (~(((((((vns_locked20 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_ready)) | (((vns_roundrobin7_grant == 2'd2) & ((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd7) & (~(((((((vns_locked23 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2)))))) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_ready));
assign soc_videooverlaysoc_videooverlaysoc_port_wdata_ready = vns_new_master_wdata_ready2;
assign soc_videooverlaysoc_litedramcrossbar_wdata_ready = vns_new_master_wdata_ready5;
assign soc_videooverlaysoc_out_dram_port_wdata_ready = vns_new_master_wdata_ready8;
assign soc_videooverlaysoc_videooverlaysoc_port_rdata_valid = vns_new_master_rdata_valid9;
assign soc_videooverlaysoc_litedramcrossbar_rdata_valid = vns_new_master_rdata_valid19;
assign soc_videooverlaysoc_out_dram_port_rdata_valid = vns_new_master_rdata_valid29;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata <= 256'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata_we <= 32'd0;
	case ({vns_new_master_wdata_ready8, vns_new_master_wdata_ready5, vns_new_master_wdata_ready2})
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata <= soc_videooverlaysoc_videooverlaysoc_port_wdata_payload_data;
			soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata_we <= soc_videooverlaysoc_videooverlaysoc_port_wdata_payload_we;
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata <= soc_videooverlaysoc_litedramcrossbar_wdata_payload_data;
			soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata_we <= soc_videooverlaysoc_litedramcrossbar_wdata_payload_we;
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata <= soc_videooverlaysoc_out_dram_port_wdata_payload_data;
			soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata_we <= soc_videooverlaysoc_out_dram_port_wdata_payload_we;
		end
		default: begin
			soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata <= 1'd0;
			soc_videooverlaysoc_videooverlaysoc_sdram_interface_wdata_we <= 1'd0;
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_port_rdata_payload_data = soc_videooverlaysoc_videooverlaysoc_sdram_interface_rdata;
assign soc_videooverlaysoc_litedramcrossbar_rdata_payload_data = soc_videooverlaysoc_videooverlaysoc_sdram_interface_rdata;
assign soc_videooverlaysoc_out_dram_port_rdata_payload_data = soc_videooverlaysoc_videooverlaysoc_sdram_interface_rdata;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_din = {soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_last, soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_first, soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_payload_addr, soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_payload_we};
assign {soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_last, soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_first, soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_payload_addr, soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_payload_we} = soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_dout;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_ready = soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_writable;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_we = soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_valid;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_first = soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_first;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_last = soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_last;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_payload_we = soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_payload_we;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_in_payload_addr = soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_payload_addr;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_source_valid = soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_readable;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_source_first = soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_first;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_source_last = soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_last;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_source_payload_we = soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_payload_we;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_source_payload_addr = soc_videooverlaysoc_out_dram_port_cmd_fifo_fifo_out_payload_addr;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_re = soc_videooverlaysoc_out_dram_port_cmd_fifo_source_ready;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_ce = (soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_writable & soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_we);
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_ce = (soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_readable & soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_re);
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_writable = (((soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q[2] == soc_videooverlaysoc_out_dram_port_cmd_fifo_consume_wdomain[2]) | (soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q[1] == soc_videooverlaysoc_out_dram_port_cmd_fifo_consume_wdomain[1])) | (soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q[0] != soc_videooverlaysoc_out_dram_port_cmd_fifo_consume_wdomain[0]));
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_readable = (soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q != soc_videooverlaysoc_out_dram_port_cmd_fifo_produce_rdomain);
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_adr = soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_binary[1:0];
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_dat_w = soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_din;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_we = soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_ce;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_rdport_adr = soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next_binary[1:0];
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_asyncfifo_dout = soc_videooverlaysoc_out_dram_port_cmd_fifo_rdport_dat_r;
always @(*) begin
	soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_next_binary <= 3'd0;
	if (soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_ce) begin
		soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_next_binary <= (soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_next_binary <= soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_binary;
	end
end
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_next = (soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_next_binary ^ soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_next_binary[2:1]);
always @(*) begin
	soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next_binary <= 3'd0;
	if (soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_ce) begin
		soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next_binary <= (soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next_binary <= soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_binary;
	end
end
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next = (soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next_binary ^ soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next_binary[2:1]);
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_valid = soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_valid;
assign soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_ready = soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_ready;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_first = soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_first;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_last = soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_last;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_payload_we = soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_payload_we;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_sink_payload_addr = soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_payload_addr;
assign soc_videooverlaysoc_out_dram_port_cmd_valid = soc_videooverlaysoc_out_dram_port_cmd_fifo_source_valid;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_source_ready = soc_videooverlaysoc_out_dram_port_cmd_ready;
assign soc_videooverlaysoc_out_dram_port_cmd_first = soc_videooverlaysoc_out_dram_port_cmd_fifo_source_first;
assign soc_videooverlaysoc_out_dram_port_cmd_last = soc_videooverlaysoc_out_dram_port_cmd_fifo_source_last;
assign soc_videooverlaysoc_out_dram_port_cmd_payload_we = soc_videooverlaysoc_out_dram_port_cmd_fifo_source_payload_we;
assign soc_videooverlaysoc_out_dram_port_cmd_payload_addr = soc_videooverlaysoc_out_dram_port_cmd_fifo_source_payload_addr;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_din = {soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_in_last, soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_in_first, soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_in_payload_data};
assign {soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_out_last, soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_out_first, soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_out_payload_data} = soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_dout;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_ready = soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_writable;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_we = soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_valid;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_in_first = soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_first;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_in_last = soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_last;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_in_payload_data = soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_payload_data;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_source_valid = soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_readable;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_source_first = soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_out_first;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_source_last = soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_out_last;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_source_payload_data = soc_videooverlaysoc_out_dram_port_rdata_fifo_fifo_out_payload_data;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_re = soc_videooverlaysoc_out_dram_port_rdata_fifo_source_ready;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_ce = (soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_writable & soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_we);
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_ce = (soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_readable & soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_re);
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_writable = (((soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q[4] == soc_videooverlaysoc_out_dram_port_rdata_fifo_consume_wdomain[4]) | (soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q[3] == soc_videooverlaysoc_out_dram_port_rdata_fifo_consume_wdomain[3])) | (soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q[2:0] != soc_videooverlaysoc_out_dram_port_rdata_fifo_consume_wdomain[2:0]));
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_readable = (soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q != soc_videooverlaysoc_out_dram_port_rdata_fifo_produce_rdomain);
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_adr = soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_binary[3:0];
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_dat_w = soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_din;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_we = soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_ce;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_rdport_adr = soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next_binary[3:0];
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_asyncfifo_dout = soc_videooverlaysoc_out_dram_port_rdata_fifo_rdport_dat_r;
always @(*) begin
	soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_next_binary <= 5'd0;
	if (soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_ce) begin
		soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_next_binary <= (soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_next_binary <= soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_binary;
	end
end
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_next = (soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_next_binary ^ soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_next_binary[4:1]);
always @(*) begin
	soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next_binary <= 5'd0;
	if (soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_ce) begin
		soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next_binary <= (soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next_binary <= soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_binary;
	end
end
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next = (soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next_binary ^ soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next_binary[4:1]);
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_valid = soc_videooverlaysoc_out_dram_port_rdata_valid;
assign soc_videooverlaysoc_out_dram_port_rdata_ready = soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_ready;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_first = soc_videooverlaysoc_out_dram_port_rdata_first;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_last = soc_videooverlaysoc_out_dram_port_rdata_last;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_sink_payload_data = soc_videooverlaysoc_out_dram_port_rdata_payload_data;
assign soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_valid = soc_videooverlaysoc_out_dram_port_rdata_fifo_source_valid;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_source_ready = soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_ready;
assign soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_first = soc_videooverlaysoc_out_dram_port_rdata_fifo_source_first;
assign soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_last = soc_videooverlaysoc_out_dram_port_rdata_fifo_source_last;
assign soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_payload_data = soc_videooverlaysoc_out_dram_port_rdata_fifo_source_payload_data;
always @(*) begin
	soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_payload_addr <= 24'd0;
	soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_ready <= 1'd0;
	soc_videooverlaysoc_out_dram_port_counter_ce <= 1'd0;
	soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_valid <= 1'd0;
	if (soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_valid) begin
		if ((soc_videooverlaysoc_out_dram_port_counter == 1'd0)) begin
			soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_valid <= 1'd1;
			soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_payload_addr <= soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_payload_addr[26:3];
			soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_ready <= soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_ready;
			soc_videooverlaysoc_out_dram_port_counter_ce <= soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_ready;
		end else begin
			soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_ready <= 1'd1;
			soc_videooverlaysoc_out_dram_port_counter_ce <= 1'd1;
		end
	end
end
always @(*) begin
	soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_valid <= 1'd0;
	soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_payload_sel <= 8'd0;
	if ((soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_valid & soc_videooverlaysoc_out_dram_port_litedramnativeport0_cmd_ready)) begin
		soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_valid <= 1'd1;
		soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_payload_sel <= 8'd255;
	end
end
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_valid = soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_valid;
assign soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_ready = soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_ready;
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_first = soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_first;
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_last = soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_last;
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_payload_data = soc_videooverlaysoc_out_dram_port_litedramnativeport0_rdata_payload_data;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_sink_valid = soc_videooverlaysoc_out_dram_port_rdata_buffer_source_valid;
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_source_ready = soc_videooverlaysoc_out_dram_port_rdata_converter_sink_ready;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_sink_first = soc_videooverlaysoc_out_dram_port_rdata_buffer_source_first;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_sink_last = soc_videooverlaysoc_out_dram_port_rdata_buffer_source_last;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_sink_payload_data = soc_videooverlaysoc_out_dram_port_rdata_buffer_source_payload_data;
assign soc_videooverlaysoc_out_dram_port_rdata_chunk_valid = ((soc_videooverlaysoc_out_dram_port_cmd_buffer_source_payload_sel & soc_videooverlaysoc_out_dram_port_rdata_chunk) != 1'd0);
always @(*) begin
	soc_videooverlaysoc_out_dram_port_rdata_converter_source_ready <= 1'd0;
	soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_valid <= 1'd0;
	soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_payload_data <= 32'd0;
	if (soc_videooverlaysoc_out_dram_port_litedramnativeport1_flush) begin
		soc_videooverlaysoc_out_dram_port_rdata_converter_source_ready <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_out_dram_port_cmd_buffer_source_valid) begin
			if (soc_videooverlaysoc_out_dram_port_rdata_chunk_valid) begin
				soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_valid <= soc_videooverlaysoc_out_dram_port_rdata_converter_source_valid;
				soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_payload_data <= soc_videooverlaysoc_out_dram_port_rdata_converter_source_payload_data;
				soc_videooverlaysoc_out_dram_port_rdata_converter_source_ready <= soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_ready;
			end else begin
				soc_videooverlaysoc_out_dram_port_rdata_converter_source_ready <= 1'd1;
			end
		end
	end
end
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_source_ready = (soc_videooverlaysoc_out_dram_port_rdata_converter_source_ready & soc_videooverlaysoc_out_dram_port_rdata_chunk[7]);
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_din = {soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_in_last, soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_in_first, soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_in_payload_sel};
assign {soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_out_last, soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_out_first, soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_out_payload_sel} = soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_dout;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_ready = soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_writable;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_we = soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_valid;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_in_first = soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_first;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_in_last = soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_last;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_in_payload_sel = soc_videooverlaysoc_out_dram_port_cmd_buffer_sink_payload_sel;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_source_valid = soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_readable;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_source_first = soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_out_first;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_source_last = soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_out_last;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_source_payload_sel = soc_videooverlaysoc_out_dram_port_cmd_buffer_fifo_out_payload_sel;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_re = soc_videooverlaysoc_out_dram_port_cmd_buffer_source_ready;
always @(*) begin
	soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_adr <= 2'd0;
	if (soc_videooverlaysoc_out_dram_port_cmd_buffer_replace) begin
		soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_adr <= (soc_videooverlaysoc_out_dram_port_cmd_buffer_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_adr <= soc_videooverlaysoc_out_dram_port_cmd_buffer_produce;
	end
end
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_dat_w = soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_din;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_we = (soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_we & (soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_writable | soc_videooverlaysoc_out_dram_port_cmd_buffer_replace));
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_do_read = (soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_readable & soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_re);
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_rdport_adr = soc_videooverlaysoc_out_dram_port_cmd_buffer_consume;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_dout = soc_videooverlaysoc_out_dram_port_cmd_buffer_rdport_dat_r;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_writable = (soc_videooverlaysoc_out_dram_port_cmd_buffer_level != 3'd4);
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_readable = (soc_videooverlaysoc_out_dram_port_cmd_buffer_level != 1'd0);
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_pipe_ce = (soc_videooverlaysoc_out_dram_port_rdata_buffer_source_ready | (~soc_videooverlaysoc_out_dram_port_rdata_buffer_valid_n));
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_ready = soc_videooverlaysoc_out_dram_port_rdata_buffer_pipe_ce;
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_source_valid = soc_videooverlaysoc_out_dram_port_rdata_buffer_valid_n;
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_busy = (1'd0 | soc_videooverlaysoc_out_dram_port_rdata_buffer_valid_n);
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_source_first = soc_videooverlaysoc_out_dram_port_rdata_buffer_first_n;
assign soc_videooverlaysoc_out_dram_port_rdata_buffer_source_last = soc_videooverlaysoc_out_dram_port_rdata_buffer_last_n;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_valid = soc_videooverlaysoc_out_dram_port_rdata_converter_sink_valid;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_first = soc_videooverlaysoc_out_dram_port_rdata_converter_sink_first;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_last = soc_videooverlaysoc_out_dram_port_rdata_converter_sink_last;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_sink_ready = soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_ready;
always @(*) begin
	soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data <= 256'd0;
	soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[31:0] <= soc_videooverlaysoc_out_dram_port_rdata_converter_sink_payload_data[31:0];
	soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[63:32] <= soc_videooverlaysoc_out_dram_port_rdata_converter_sink_payload_data[63:32];
	soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[95:64] <= soc_videooverlaysoc_out_dram_port_rdata_converter_sink_payload_data[95:64];
	soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[127:96] <= soc_videooverlaysoc_out_dram_port_rdata_converter_sink_payload_data[127:96];
	soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[159:128] <= soc_videooverlaysoc_out_dram_port_rdata_converter_sink_payload_data[159:128];
	soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[191:160] <= soc_videooverlaysoc_out_dram_port_rdata_converter_sink_payload_data[191:160];
	soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[223:192] <= soc_videooverlaysoc_out_dram_port_rdata_converter_sink_payload_data[223:192];
	soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[255:224] <= soc_videooverlaysoc_out_dram_port_rdata_converter_sink_payload_data[255:224];
end
assign soc_videooverlaysoc_out_dram_port_rdata_converter_source_valid = soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_valid;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_source_first = soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_first;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_source_last = soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_last;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_ready = soc_videooverlaysoc_out_dram_port_rdata_converter_source_ready;
assign {soc_videooverlaysoc_out_dram_port_rdata_converter_source_payload_data} = soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_payload_data;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_valid = soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_valid;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_ready = soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_ready;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_first = soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_first;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_last = soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_last;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_source_source_payload_data = soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_first = (soc_videooverlaysoc_out_dram_port_rdata_converter_converter_mux == 1'd0);
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_last = (soc_videooverlaysoc_out_dram_port_rdata_converter_converter_mux == 3'd7);
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_valid = soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_valid;
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_first = (soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_first & soc_videooverlaysoc_out_dram_port_rdata_converter_converter_first);
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_last = (soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_last & soc_videooverlaysoc_out_dram_port_rdata_converter_converter_last);
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_ready = (soc_videooverlaysoc_out_dram_port_rdata_converter_converter_last & soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_ready);
always @(*) begin
	soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data <= 32'd0;
	case (soc_videooverlaysoc_out_dram_port_rdata_converter_converter_mux)
		1'd0: begin
			soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data <= soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[255:224];
		end
		1'd1: begin
			soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data <= soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[223:192];
		end
		2'd2: begin
			soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data <= soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[191:160];
		end
		2'd3: begin
			soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data <= soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[159:128];
		end
		3'd4: begin
			soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data <= soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[127:96];
		end
		3'd5: begin
			soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data <= soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[95:64];
		end
		3'd6: begin
			soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data <= soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[63:32];
		end
		default: begin
			soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_data <= soc_videooverlaysoc_out_dram_port_rdata_converter_converter_sink_payload_data[31:0];
		end
	endcase
end
assign soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_payload_valid_token_count = soc_videooverlaysoc_out_dram_port_rdata_converter_converter_last;
assign soc_videooverlaysoc_videooverlaysoc_data_port_adr = soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[10:3];
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_data_port_dat_w <= 256'd0;
	soc_videooverlaysoc_videooverlaysoc_data_port_we <= 32'd0;
	if (soc_videooverlaysoc_videooverlaysoc_write_from_slave) begin
		soc_videooverlaysoc_videooverlaysoc_data_port_dat_w <= soc_videooverlaysoc_videooverlaysoc_dat_r;
		soc_videooverlaysoc_videooverlaysoc_data_port_we <= {32{1'd1}};
	end else begin
		soc_videooverlaysoc_videooverlaysoc_data_port_dat_w <= {8{soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_w}};
		if ((((soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_cyc & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_stb) & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_we) & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_ack)) begin
			soc_videooverlaysoc_videooverlaysoc_data_port_we <= {({4{(soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[2:0] == 1'd0)}} & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_sel), ({4{(soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[2:0] == 1'd1)}} & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_sel), ({4{(soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[2:0] == 2'd2)}} & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_sel), ({4{(soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[2:0] == 2'd3)}} & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_sel), ({4{(soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[2:0] == 3'd4)}} & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_sel), ({4{(soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[2:0] == 3'd5)}} & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_sel), ({4{(soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[2:0] == 3'd6)}} & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_sel), ({4{(soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[2:0] == 3'd7)}} & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_sel)};
		end
	end
end
assign soc_videooverlaysoc_videooverlaysoc_dat_w = soc_videooverlaysoc_videooverlaysoc_data_port_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_sel = 32'd4294967295;
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r <= 32'd0;
	case (soc_videooverlaysoc_videooverlaysoc_adr_offset_r)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[255:224];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[223:192];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[191:160];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[159:128];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[127:96];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[95:64];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[63:32];
		end
		default: begin
			soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[31:0];
		end
	endcase
end
assign {soc_videooverlaysoc_videooverlaysoc_tag_do_dirty, soc_videooverlaysoc_videooverlaysoc_tag_do_tag} = soc_videooverlaysoc_videooverlaysoc_tag_port_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_tag_port_dat_w = {soc_videooverlaysoc_videooverlaysoc_tag_di_dirty, soc_videooverlaysoc_videooverlaysoc_tag_di_tag};
assign soc_videooverlaysoc_videooverlaysoc_tag_port_adr = soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[10:3];
assign soc_videooverlaysoc_videooverlaysoc_tag_di_tag = soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[29:11];
assign soc_videooverlaysoc_videooverlaysoc_adr = {soc_videooverlaysoc_videooverlaysoc_tag_do_tag, soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[10:3]};
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_tag_di_dirty <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_word_clr <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_word_inc <= 1'd0;
	vns_fullmemorywe_next_state <= 3'd0;
	soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_ack <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_write_from_slave <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_tag_port_we <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_cyc <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_stb <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_we <= 1'd0;
	vns_fullmemorywe_next_state <= vns_fullmemorywe_state;
	case (vns_fullmemorywe_state)
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_word_clr <= 1'd1;
			if ((soc_videooverlaysoc_videooverlaysoc_tag_do_tag == soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[29:11])) begin
				soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_ack <= 1'd1;
				if (soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_we) begin
					soc_videooverlaysoc_videooverlaysoc_tag_di_dirty <= 1'd1;
					soc_videooverlaysoc_videooverlaysoc_tag_port_we <= 1'd1;
				end
				vns_fullmemorywe_next_state <= 1'd0;
			end else begin
				if (soc_videooverlaysoc_videooverlaysoc_tag_do_dirty) begin
					vns_fullmemorywe_next_state <= 2'd2;
				end else begin
					vns_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_stb <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_cyc <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_we <= 1'd1;
			if (soc_videooverlaysoc_videooverlaysoc_ack) begin
				soc_videooverlaysoc_videooverlaysoc_word_inc <= 1'd1;
				if (1'd1) begin
					vns_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_tag_port_we <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_word_clr <= 1'd1;
			vns_fullmemorywe_next_state <= 3'd4;
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_stb <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_cyc <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_we <= 1'd0;
			if (soc_videooverlaysoc_videooverlaysoc_ack) begin
				soc_videooverlaysoc_videooverlaysoc_write_from_slave <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_word_inc <= 1'd1;
				if (1'd1) begin
					vns_fullmemorywe_next_state <= 1'd1;
				end else begin
					vns_fullmemorywe_next_state <= 3'd4;
				end
			end
		end
		default: begin
			if ((soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_cyc & soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_stb)) begin
				vns_fullmemorywe_next_state <= 1'd1;
			end
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_port_wdata_payload_data <= 256'd0;
	vns_litedramwishbone2native_next_state <= 2'd0;
	soc_videooverlaysoc_videooverlaysoc_port_wdata_payload_we <= 32'd0;
	soc_videooverlaysoc_videooverlaysoc_port_rdata_ready <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_port_cmd_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_dat_r <= 256'd0;
	soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr <= 24'd0;
	soc_videooverlaysoc_videooverlaysoc_port_wdata_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_ack <= 1'd0;
	vns_litedramwishbone2native_next_state <= vns_litedramwishbone2native_state;
	case (vns_litedramwishbone2native_state)
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_port_cmd_valid <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr <= soc_videooverlaysoc_videooverlaysoc_adr;
			soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we <= soc_videooverlaysoc_videooverlaysoc_we;
			if (soc_videooverlaysoc_videooverlaysoc_port_cmd_ready) begin
				if (soc_videooverlaysoc_videooverlaysoc_we) begin
					vns_litedramwishbone2native_next_state <= 2'd2;
				end else begin
					vns_litedramwishbone2native_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_port_wdata_valid <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_port_wdata_payload_we <= soc_videooverlaysoc_videooverlaysoc_sel;
			soc_videooverlaysoc_videooverlaysoc_port_wdata_payload_data <= soc_videooverlaysoc_videooverlaysoc_dat_w;
			if (soc_videooverlaysoc_videooverlaysoc_port_wdata_ready) begin
				soc_videooverlaysoc_videooverlaysoc_ack <= 1'd1;
				vns_litedramwishbone2native_next_state <= 1'd0;
			end
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_port_rdata_ready <= 1'd1;
			if (soc_videooverlaysoc_videooverlaysoc_port_rdata_valid) begin
				soc_videooverlaysoc_videooverlaysoc_dat_r <= soc_videooverlaysoc_videooverlaysoc_port_rdata_payload_data;
				soc_videooverlaysoc_videooverlaysoc_ack <= 1'd1;
				vns_litedramwishbone2native_next_state <= 1'd0;
			end
		end
		default: begin
			if ((soc_videooverlaysoc_videooverlaysoc_cyc & soc_videooverlaysoc_videooverlaysoc_stb)) begin
				vns_litedramwishbone2native_next_state <= 1'd1;
			end
		end
	endcase
end
assign hdmi_in0_freq_fmeter_clk = soc_videooverlaysoc_hdmi_in0_freq_clk0;
assign soc_videooverlaysoc_hdmi_in0_freq_period_done = (soc_videooverlaysoc_hdmi_in0_freq_period_counter == 27'd100000000);
assign soc_videooverlaysoc_hdmi_in0_freq_ce = 1'd1;
assign soc_videooverlaysoc_hdmi_in0_freq_sampler_latch = soc_videooverlaysoc_hdmi_in0_freq_period_done;
assign soc_videooverlaysoc_hdmi_in0_freq_sampler_i = soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o;
assign soc_videooverlaysoc_hdmi_in0_freq_status = soc_videooverlaysoc_hdmi_in0_freq_sampler_o;
always @(*) begin
	soc_videooverlaysoc_hdmi_in0_freq_q_next_binary <= 6'd0;
	if (soc_videooverlaysoc_hdmi_in0_freq_ce) begin
		soc_videooverlaysoc_hdmi_in0_freq_q_next_binary <= (soc_videooverlaysoc_hdmi_in0_freq_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_hdmi_in0_freq_q_next_binary <= soc_videooverlaysoc_hdmi_in0_freq_q_binary;
	end
end
assign soc_videooverlaysoc_hdmi_in0_freq_q_next = (soc_videooverlaysoc_hdmi_in0_freq_q_next_binary ^ soc_videooverlaysoc_hdmi_in0_freq_q_next_binary[5:1]);
always @(*) begin
	soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb <= 6'd0;
	soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[5] <= soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_i[5];
	soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[4] <= (soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[5] ^ soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_i[4]);
	soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[3] <= (soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[4] ^ soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_i[3]);
	soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[2] <= (soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[3] ^ soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_i[2]);
	soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[1] <= (soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[2] ^ soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_i[1]);
	soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[0] <= (soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb[1] ^ soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_i[0]);
end
assign soc_videooverlaysoc_hdmi_in0_freq_sampler_inc = (soc_videooverlaysoc_hdmi_in0_freq_sampler_i - soc_videooverlaysoc_hdmi_in0_freq_sampler_i_d);
assign soc_videooverlaysoc_hdmi_in0_charsync0_raw_data = soc_videooverlaysoc_hdmi_in0_s7datacapture0_d;
assign soc_videooverlaysoc_hdmi_in0_wer0_data = soc_videooverlaysoc_hdmi_in0_charsync0_data;
assign soc_videooverlaysoc_hdmi_in0_decoding0_valid_i = soc_videooverlaysoc_hdmi_in0_charsync0_synced;
assign soc_videooverlaysoc_hdmi_in0_decoding0_input = soc_videooverlaysoc_hdmi_in0_charsync0_data;
assign soc_videooverlaysoc_hdmi_in0_charsync1_raw_data = soc_videooverlaysoc_hdmi_in0_s7datacapture1_d;
assign soc_videooverlaysoc_hdmi_in0_wer1_data = soc_videooverlaysoc_hdmi_in0_charsync1_data;
assign soc_videooverlaysoc_hdmi_in0_decoding1_valid_i = soc_videooverlaysoc_hdmi_in0_charsync1_synced;
assign soc_videooverlaysoc_hdmi_in0_decoding1_input = soc_videooverlaysoc_hdmi_in0_charsync1_data;
assign soc_videooverlaysoc_hdmi_in0_charsync2_raw_data = soc_videooverlaysoc_hdmi_in0_s7datacapture2_d;
assign soc_videooverlaysoc_hdmi_in0_wer2_data = soc_videooverlaysoc_hdmi_in0_charsync2_data;
assign soc_videooverlaysoc_hdmi_in0_decoding2_valid_i = soc_videooverlaysoc_hdmi_in0_charsync2_synced;
assign soc_videooverlaysoc_hdmi_in0_decoding2_input = soc_videooverlaysoc_hdmi_in0_charsync2_data;
assign soc_videooverlaysoc_hdmi_in0_chansync_valid_i = ((soc_videooverlaysoc_hdmi_in0_decoding0_valid_o & soc_videooverlaysoc_hdmi_in0_decoding1_valid_o) & soc_videooverlaysoc_hdmi_in0_decoding2_valid_o);
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in0_raw = soc_videooverlaysoc_hdmi_in0_decoding0_output_raw;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in0_d = soc_videooverlaysoc_hdmi_in0_decoding0_output_d;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in0_c = soc_videooverlaysoc_hdmi_in0_decoding0_output_c;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in0_de = soc_videooverlaysoc_hdmi_in0_decoding0_output_de;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in1_raw = soc_videooverlaysoc_hdmi_in0_decoding1_output_raw;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in1_d = soc_videooverlaysoc_hdmi_in0_decoding1_output_d;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in1_c = soc_videooverlaysoc_hdmi_in0_decoding1_output_c;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in1_de = soc_videooverlaysoc_hdmi_in0_decoding1_output_de;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in2_raw = soc_videooverlaysoc_hdmi_in0_decoding2_output_raw;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in2_d = soc_videooverlaysoc_hdmi_in0_decoding2_output_d;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in2_c = soc_videooverlaysoc_hdmi_in0_decoding2_output_c;
assign soc_videooverlaysoc_hdmi_in0_chansync_data_in2_de = soc_videooverlaysoc_hdmi_in0_decoding2_output_de;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_valid_i = soc_videooverlaysoc_hdmi_in0_chansync_chan_synced;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_raw = soc_videooverlaysoc_hdmi_in0_chansync_data_out0_raw;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_d = soc_videooverlaysoc_hdmi_in0_chansync_data_out0_d;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_c = soc_videooverlaysoc_hdmi_in0_chansync_data_out0_c;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_de = soc_videooverlaysoc_hdmi_in0_chansync_data_out0_de;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_raw = soc_videooverlaysoc_hdmi_in0_chansync_data_out1_raw;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_d = soc_videooverlaysoc_hdmi_in0_chansync_data_out1_d;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_c = soc_videooverlaysoc_hdmi_in0_chansync_data_out1_c;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_de = soc_videooverlaysoc_hdmi_in0_chansync_data_out1_de;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_raw = soc_videooverlaysoc_hdmi_in0_chansync_data_out2_raw;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_d = soc_videooverlaysoc_hdmi_in0_chansync_data_out2_d;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_c = soc_videooverlaysoc_hdmi_in0_chansync_data_out2_c;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_de = soc_videooverlaysoc_hdmi_in0_chansync_data_out2_de;
assign soc_videooverlaysoc_hdmi_in0_syncpol_de_int = soc_videooverlaysoc_hdmi_in0_decode_terc4_de_o;
assign soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_raw = soc_videooverlaysoc_hdmi_in0_chansync_data_out0_raw;
assign soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_d = soc_videooverlaysoc_hdmi_in0_chansync_data_out0_d;
assign soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_c = soc_videooverlaysoc_hdmi_in0_chansync_data_out0_c;
assign soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_de = soc_videooverlaysoc_hdmi_in0_chansync_data_out0_de;
assign soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_raw = soc_videooverlaysoc_hdmi_in0_chansync_data_out1_raw;
assign soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_d = soc_videooverlaysoc_hdmi_in0_chansync_data_out1_d;
assign soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_c = soc_videooverlaysoc_hdmi_in0_chansync_data_out1_c;
assign soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_de = soc_videooverlaysoc_hdmi_in0_chansync_data_out1_de;
assign soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_raw = soc_videooverlaysoc_hdmi_in0_chansync_data_out2_raw;
assign soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_d = soc_videooverlaysoc_hdmi_in0_chansync_data_out2_d;
assign soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_c = soc_videooverlaysoc_hdmi_in0_chansync_data_out2_c;
assign soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_de = soc_videooverlaysoc_hdmi_in0_chansync_data_out2_de;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_raw = soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_raw;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_d = soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_d;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_c = soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_c;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_de = soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_de;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in1_raw = soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_raw;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in1_d = soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_d;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in1_c = soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_c;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in1_de = soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_de;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in2_raw = soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_raw;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in2_d = soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_d;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in2_c = soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_c;
assign soc_videooverlaysoc_hdmi_in0_syncpol_data_in2_de = soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_de;
assign soc_videooverlaysoc_hdmi_in0_syncpol_valid_i = soc_videooverlaysoc_hdmi_in0_chansync_chan_synced;
assign soc_videooverlaysoc_hdmi_in0_resdetection_valid_i = soc_videooverlaysoc_hdmi_in0_syncpol_valid_o;
assign soc_videooverlaysoc_hdmi_in0_resdetection_de = soc_videooverlaysoc_hdmi_in0_syncpol_de;
assign soc_videooverlaysoc_hdmi_in0_resdetection_vsync = soc_videooverlaysoc_hdmi_in0_syncpol_vsync;
assign soc_videooverlaysoc_hdmi_in0_edid_hpd_notif_n = (~hdmi_in0_hpd_notif);
assign soc_videooverlaysoc_hdmi_in0_edid_sda_o = (~soc_videooverlaysoc_hdmi_in0_edid_sda_drv_reg);
assign soc_videooverlaysoc_hdmi_in0_edid_scl_rising = (soc_videooverlaysoc_hdmi_in0_edid_scl_i & (~soc_videooverlaysoc_hdmi_in0_edid_scl_r));
assign soc_videooverlaysoc_hdmi_in0_edid_sda_rising = (soc_videooverlaysoc_hdmi_in0_edid_sda_i & (~soc_videooverlaysoc_hdmi_in0_edid_sda_r));
assign soc_videooverlaysoc_hdmi_in0_edid_sda_falling = ((~soc_videooverlaysoc_hdmi_in0_edid_sda_i) & soc_videooverlaysoc_hdmi_in0_edid_sda_r);
assign soc_videooverlaysoc_hdmi_in0_edid_start = (soc_videooverlaysoc_hdmi_in0_edid_scl_i & soc_videooverlaysoc_hdmi_in0_edid_sda_falling);
assign soc_videooverlaysoc_hdmi_in0_edid_adr = soc_videooverlaysoc_hdmi_in0_edid_offset_counter;
always @(*) begin
	soc_videooverlaysoc_hdmi_in0_edid_sda_drv <= 1'd0;
	if (soc_videooverlaysoc_hdmi_in0_edid_zero_drv) begin
		soc_videooverlaysoc_hdmi_in0_edid_sda_drv <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_hdmi_in0_edid_data_drv) begin
			soc_videooverlaysoc_hdmi_in0_edid_sda_drv <= (~soc_videooverlaysoc_hdmi_in0_edid_data_bit);
		end
	end
end
always @(*) begin
	soc_videooverlaysoc_hdmi_in0_edid_update_is_read <= 1'd0;
	vns_edid0_next_state <= 4'd0;
	soc_videooverlaysoc_hdmi_in0_edid_zero_drv <= 1'd0;
	soc_videooverlaysoc_hdmi_in0_edid_oc_load <= 1'd0;
	soc_videooverlaysoc_hdmi_in0_edid_oc_inc <= 1'd0;
	soc_videooverlaysoc_hdmi_in0_edid_data_drv_en <= 1'd0;
	soc_videooverlaysoc_hdmi_in0_edid_data_drv_stop <= 1'd0;
	vns_edid0_next_state <= vns_edid0_state;
	case (vns_edid0_state)
		1'd1: begin
			if ((soc_videooverlaysoc_hdmi_in0_edid_counter == 4'd8)) begin
				if ((soc_videooverlaysoc_hdmi_in0_edid_din[7:1] == 7'd80)) begin
					soc_videooverlaysoc_hdmi_in0_edid_update_is_read <= 1'd1;
					vns_edid0_next_state <= 2'd2;
				end else begin
					vns_edid0_next_state <= 1'd0;
				end
			end
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
		2'd2: begin
			if ((~soc_videooverlaysoc_hdmi_in0_edid_scl_i)) begin
				vns_edid0_next_state <= 2'd3;
			end
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in0_edid_zero_drv <= 1'd1;
			if (soc_videooverlaysoc_hdmi_in0_edid_scl_i) begin
				vns_edid0_next_state <= 3'd4;
			end
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in0_edid_zero_drv <= 1'd1;
			if ((~soc_videooverlaysoc_hdmi_in0_edid_scl_i)) begin
				if (soc_videooverlaysoc_hdmi_in0_edid_is_read) begin
					vns_edid0_next_state <= 4'd9;
				end else begin
					vns_edid0_next_state <= 3'd5;
				end
			end
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
		3'd5: begin
			if ((soc_videooverlaysoc_hdmi_in0_edid_counter == 4'd8)) begin
				soc_videooverlaysoc_hdmi_in0_edid_oc_load <= 1'd1;
				vns_edid0_next_state <= 3'd6;
			end
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
		3'd6: begin
			if ((~soc_videooverlaysoc_hdmi_in0_edid_scl_i)) begin
				vns_edid0_next_state <= 3'd7;
			end
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in0_edid_zero_drv <= 1'd1;
			if (soc_videooverlaysoc_hdmi_in0_edid_scl_i) begin
				vns_edid0_next_state <= 4'd8;
			end
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
		4'd8: begin
			soc_videooverlaysoc_hdmi_in0_edid_zero_drv <= 1'd1;
			if ((~soc_videooverlaysoc_hdmi_in0_edid_scl_i)) begin
				vns_edid0_next_state <= 1'd1;
			end
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
		4'd9: begin
			if ((~soc_videooverlaysoc_hdmi_in0_edid_scl_i)) begin
				if ((soc_videooverlaysoc_hdmi_in0_edid_counter == 4'd8)) begin
					soc_videooverlaysoc_hdmi_in0_edid_data_drv_stop <= 1'd1;
					vns_edid0_next_state <= 4'd10;
				end else begin
					soc_videooverlaysoc_hdmi_in0_edid_data_drv_en <= 1'd1;
				end
			end
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
		4'd10: begin
			if (soc_videooverlaysoc_hdmi_in0_edid_scl_rising) begin
				soc_videooverlaysoc_hdmi_in0_edid_oc_inc <= 1'd1;
				if (soc_videooverlaysoc_hdmi_in0_edid_sda_i) begin
					vns_edid0_next_state <= 1'd0;
				end else begin
					vns_edid0_next_state <= 4'd9;
				end
			end
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
		default: begin
			if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
				vns_edid0_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_hdmi_in0_locked_status = soc_videooverlaysoc_hdmi_in0_locked;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_d = (~soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_q);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_d = soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_q;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i = soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_d = soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_mdata = soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_sdata = soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_d;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_too_late = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_lateness == 8'd255);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_too_early = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_lateness == 1'd0);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_rst = soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_master_inc = soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_master_ce = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_o | soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_o);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_slave_inc = soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_slave_ce = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_o | soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_o);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_r[0]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_r[1]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_r[2]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_r[3]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_r[4]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_reset_lateness = soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_i = soc_videooverlaysoc_hdmi_in0_s7datacapture0_phase_reset_re;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst = (hdmi_in0_pix1p25x_rst | hdmi_in0_pix_rst);
assign hdmi_in0_data0_cap_write_clk = hdmi_in0_pix1p25x_clk;
assign hdmi_in0_data0_cap_read_clk = hdmi_in0_pix_clk;
assign hdmi_in0_data0_cap_write_rst = soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst_write;
assign hdmi_in0_data0_cap_read_rst = soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst_read;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_transition = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_mdata_d != soc_videooverlaysoc_hdmi_in0_s7datacapture0_mdata);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_inc = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_transition & (soc_videooverlaysoc_hdmi_in0_s7datacapture0_mdata == soc_videooverlaysoc_hdmi_in0_s7datacapture0_sdata));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_dec = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_transition & (soc_videooverlaysoc_hdmi_in0_s7datacapture0_mdata != soc_videooverlaysoc_hdmi_in0_s7datacapture0_sdata));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_charsync0_raw = {soc_videooverlaysoc_hdmi_in0_charsync0_raw_data, soc_videooverlaysoc_hdmi_in0_charsync0_raw_data1};
always @(*) begin
	soc_videooverlaysoc_hdmi_in0_wer0_transitions <= 8'd0;
	soc_videooverlaysoc_hdmi_in0_wer0_transitions[0] <= (soc_videooverlaysoc_hdmi_in0_wer0_data_r[0] ^ soc_videooverlaysoc_hdmi_in0_wer0_data_r[1]);
	soc_videooverlaysoc_hdmi_in0_wer0_transitions[1] <= (soc_videooverlaysoc_hdmi_in0_wer0_data_r[1] ^ soc_videooverlaysoc_hdmi_in0_wer0_data_r[2]);
	soc_videooverlaysoc_hdmi_in0_wer0_transitions[2] <= (soc_videooverlaysoc_hdmi_in0_wer0_data_r[2] ^ soc_videooverlaysoc_hdmi_in0_wer0_data_r[3]);
	soc_videooverlaysoc_hdmi_in0_wer0_transitions[3] <= (soc_videooverlaysoc_hdmi_in0_wer0_data_r[3] ^ soc_videooverlaysoc_hdmi_in0_wer0_data_r[4]);
	soc_videooverlaysoc_hdmi_in0_wer0_transitions[4] <= (soc_videooverlaysoc_hdmi_in0_wer0_data_r[4] ^ soc_videooverlaysoc_hdmi_in0_wer0_data_r[5]);
	soc_videooverlaysoc_hdmi_in0_wer0_transitions[5] <= (soc_videooverlaysoc_hdmi_in0_wer0_data_r[5] ^ soc_videooverlaysoc_hdmi_in0_wer0_data_r[6]);
	soc_videooverlaysoc_hdmi_in0_wer0_transitions[6] <= (soc_videooverlaysoc_hdmi_in0_wer0_data_r[6] ^ soc_videooverlaysoc_hdmi_in0_wer0_data_r[7]);
	soc_videooverlaysoc_hdmi_in0_wer0_transitions[7] <= (soc_videooverlaysoc_hdmi_in0_wer0_data_r[7] ^ soc_videooverlaysoc_hdmi_in0_wer0_data_r[8]);
end
assign soc_videooverlaysoc_hdmi_in0_wer0_i = soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_r_updated;
assign soc_videooverlaysoc_hdmi_in0_wer0_o = (soc_videooverlaysoc_hdmi_in0_wer0_toggle_o ^ soc_videooverlaysoc_hdmi_in0_wer0_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_d = (~soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_q);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_d = soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_q;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i = soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_d = soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_mdata = soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_sdata = soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_d;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_too_late = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_lateness == 8'd255);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_too_early = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_lateness == 1'd0);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_rst = soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_master_inc = soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_master_ce = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_o | soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_o);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_slave_inc = soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_slave_ce = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_o | soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_o);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_r[0]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_r[1]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_r[2]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_r[3]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_r[4]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_reset_lateness = soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_i = soc_videooverlaysoc_hdmi_in0_s7datacapture1_phase_reset_re;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst = (hdmi_in0_pix1p25x_rst | hdmi_in0_pix_rst);
assign hdmi_in0_data1_cap_write_clk = hdmi_in0_pix1p25x_clk;
assign hdmi_in0_data1_cap_read_clk = hdmi_in0_pix_clk;
assign hdmi_in0_data1_cap_write_rst = soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst_write;
assign hdmi_in0_data1_cap_read_rst = soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst_read;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_transition = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_mdata_d != soc_videooverlaysoc_hdmi_in0_s7datacapture1_mdata);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_inc = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_transition & (soc_videooverlaysoc_hdmi_in0_s7datacapture1_mdata == soc_videooverlaysoc_hdmi_in0_s7datacapture1_sdata));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_dec = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_transition & (soc_videooverlaysoc_hdmi_in0_s7datacapture1_mdata != soc_videooverlaysoc_hdmi_in0_s7datacapture1_sdata));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_charsync1_raw = {soc_videooverlaysoc_hdmi_in0_charsync1_raw_data, soc_videooverlaysoc_hdmi_in0_charsync1_raw_data1};
always @(*) begin
	soc_videooverlaysoc_hdmi_in0_wer1_transitions <= 8'd0;
	soc_videooverlaysoc_hdmi_in0_wer1_transitions[0] <= (soc_videooverlaysoc_hdmi_in0_wer1_data_r[0] ^ soc_videooverlaysoc_hdmi_in0_wer1_data_r[1]);
	soc_videooverlaysoc_hdmi_in0_wer1_transitions[1] <= (soc_videooverlaysoc_hdmi_in0_wer1_data_r[1] ^ soc_videooverlaysoc_hdmi_in0_wer1_data_r[2]);
	soc_videooverlaysoc_hdmi_in0_wer1_transitions[2] <= (soc_videooverlaysoc_hdmi_in0_wer1_data_r[2] ^ soc_videooverlaysoc_hdmi_in0_wer1_data_r[3]);
	soc_videooverlaysoc_hdmi_in0_wer1_transitions[3] <= (soc_videooverlaysoc_hdmi_in0_wer1_data_r[3] ^ soc_videooverlaysoc_hdmi_in0_wer1_data_r[4]);
	soc_videooverlaysoc_hdmi_in0_wer1_transitions[4] <= (soc_videooverlaysoc_hdmi_in0_wer1_data_r[4] ^ soc_videooverlaysoc_hdmi_in0_wer1_data_r[5]);
	soc_videooverlaysoc_hdmi_in0_wer1_transitions[5] <= (soc_videooverlaysoc_hdmi_in0_wer1_data_r[5] ^ soc_videooverlaysoc_hdmi_in0_wer1_data_r[6]);
	soc_videooverlaysoc_hdmi_in0_wer1_transitions[6] <= (soc_videooverlaysoc_hdmi_in0_wer1_data_r[6] ^ soc_videooverlaysoc_hdmi_in0_wer1_data_r[7]);
	soc_videooverlaysoc_hdmi_in0_wer1_transitions[7] <= (soc_videooverlaysoc_hdmi_in0_wer1_data_r[7] ^ soc_videooverlaysoc_hdmi_in0_wer1_data_r[8]);
end
assign soc_videooverlaysoc_hdmi_in0_wer1_i = soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_r_updated;
assign soc_videooverlaysoc_hdmi_in0_wer1_o = (soc_videooverlaysoc_hdmi_in0_wer1_toggle_o ^ soc_videooverlaysoc_hdmi_in0_wer1_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_d = (~soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_q);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_d = soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_q;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i = soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_d = soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_mdata = soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_sdata = soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_d;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_too_late = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_lateness == 8'd255);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_too_early = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_lateness == 1'd0);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_rst = soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_master_inc = soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_master_ce = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_o | soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_o);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_slave_inc = soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_slave_ce = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_o | soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_o);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_r[0]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_r[1]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_r[2]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_r[3]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_i = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_re & soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_r[4]);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_reset_lateness = soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_o;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_i = soc_videooverlaysoc_hdmi_in0_s7datacapture2_phase_reset_re;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst = (hdmi_in0_pix1p25x_rst | hdmi_in0_pix_rst);
assign hdmi_in0_data2_cap_write_clk = hdmi_in0_pix1p25x_clk;
assign hdmi_in0_data2_cap_read_clk = hdmi_in0_pix_clk;
assign hdmi_in0_data2_cap_write_rst = soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst_write;
assign hdmi_in0_data2_cap_read_rst = soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst_read;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_transition = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_mdata_d != soc_videooverlaysoc_hdmi_in0_s7datacapture2_mdata);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_inc = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_transition & (soc_videooverlaysoc_hdmi_in0_s7datacapture2_mdata == soc_videooverlaysoc_hdmi_in0_s7datacapture2_sdata));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_dec = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_transition & (soc_videooverlaysoc_hdmi_in0_s7datacapture2_mdata != soc_videooverlaysoc_hdmi_in0_s7datacapture2_sdata));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_o = (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_o ^ soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_charsync2_raw = {soc_videooverlaysoc_hdmi_in0_charsync2_raw_data, soc_videooverlaysoc_hdmi_in0_charsync2_raw_data1};
always @(*) begin
	soc_videooverlaysoc_hdmi_in0_wer2_transitions <= 8'd0;
	soc_videooverlaysoc_hdmi_in0_wer2_transitions[0] <= (soc_videooverlaysoc_hdmi_in0_wer2_data_r[0] ^ soc_videooverlaysoc_hdmi_in0_wer2_data_r[1]);
	soc_videooverlaysoc_hdmi_in0_wer2_transitions[1] <= (soc_videooverlaysoc_hdmi_in0_wer2_data_r[1] ^ soc_videooverlaysoc_hdmi_in0_wer2_data_r[2]);
	soc_videooverlaysoc_hdmi_in0_wer2_transitions[2] <= (soc_videooverlaysoc_hdmi_in0_wer2_data_r[2] ^ soc_videooverlaysoc_hdmi_in0_wer2_data_r[3]);
	soc_videooverlaysoc_hdmi_in0_wer2_transitions[3] <= (soc_videooverlaysoc_hdmi_in0_wer2_data_r[3] ^ soc_videooverlaysoc_hdmi_in0_wer2_data_r[4]);
	soc_videooverlaysoc_hdmi_in0_wer2_transitions[4] <= (soc_videooverlaysoc_hdmi_in0_wer2_data_r[4] ^ soc_videooverlaysoc_hdmi_in0_wer2_data_r[5]);
	soc_videooverlaysoc_hdmi_in0_wer2_transitions[5] <= (soc_videooverlaysoc_hdmi_in0_wer2_data_r[5] ^ soc_videooverlaysoc_hdmi_in0_wer2_data_r[6]);
	soc_videooverlaysoc_hdmi_in0_wer2_transitions[6] <= (soc_videooverlaysoc_hdmi_in0_wer2_data_r[6] ^ soc_videooverlaysoc_hdmi_in0_wer2_data_r[7]);
	soc_videooverlaysoc_hdmi_in0_wer2_transitions[7] <= (soc_videooverlaysoc_hdmi_in0_wer2_data_r[7] ^ soc_videooverlaysoc_hdmi_in0_wer2_data_r[8]);
end
assign soc_videooverlaysoc_hdmi_in0_wer2_i = soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_r_updated;
assign soc_videooverlaysoc_hdmi_in0_wer2_o = (soc_videooverlaysoc_hdmi_in0_wer2_toggle_o ^ soc_videooverlaysoc_hdmi_in0_wer2_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_din = {soc_videooverlaysoc_hdmi_in0_chansync_data_in0_de, soc_videooverlaysoc_hdmi_in0_chansync_data_in0_c, soc_videooverlaysoc_hdmi_in0_chansync_data_in0_d, soc_videooverlaysoc_hdmi_in0_chansync_data_in0_raw};
assign {soc_videooverlaysoc_hdmi_in0_chansync_data_out0_de, soc_videooverlaysoc_hdmi_in0_chansync_data_out0_c, soc_videooverlaysoc_hdmi_in0_chansync_data_out0_d, soc_videooverlaysoc_hdmi_in0_chansync_data_out0_raw} = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_dout;
assign soc_videooverlaysoc_hdmi_in0_chansync_is_control0 = (~soc_videooverlaysoc_hdmi_in0_chansync_data_out0_de);
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_re = ((~soc_videooverlaysoc_hdmi_in0_chansync_is_control0) | soc_videooverlaysoc_hdmi_in0_chansync_all_control);
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_din = {soc_videooverlaysoc_hdmi_in0_chansync_data_in1_de, soc_videooverlaysoc_hdmi_in0_chansync_data_in1_c, soc_videooverlaysoc_hdmi_in0_chansync_data_in1_d, soc_videooverlaysoc_hdmi_in0_chansync_data_in1_raw};
assign {soc_videooverlaysoc_hdmi_in0_chansync_data_out1_de, soc_videooverlaysoc_hdmi_in0_chansync_data_out1_c, soc_videooverlaysoc_hdmi_in0_chansync_data_out1_d, soc_videooverlaysoc_hdmi_in0_chansync_data_out1_raw} = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_dout;
assign soc_videooverlaysoc_hdmi_in0_chansync_is_control1 = (~soc_videooverlaysoc_hdmi_in0_chansync_data_out1_de);
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_re = ((~soc_videooverlaysoc_hdmi_in0_chansync_is_control1) | soc_videooverlaysoc_hdmi_in0_chansync_all_control);
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_din = {soc_videooverlaysoc_hdmi_in0_chansync_data_in2_de, soc_videooverlaysoc_hdmi_in0_chansync_data_in2_c, soc_videooverlaysoc_hdmi_in0_chansync_data_in2_d, soc_videooverlaysoc_hdmi_in0_chansync_data_in2_raw};
assign {soc_videooverlaysoc_hdmi_in0_chansync_data_out2_de, soc_videooverlaysoc_hdmi_in0_chansync_data_out2_c, soc_videooverlaysoc_hdmi_in0_chansync_data_out2_d, soc_videooverlaysoc_hdmi_in0_chansync_data_out2_raw} = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_dout;
assign soc_videooverlaysoc_hdmi_in0_chansync_is_control2 = (~soc_videooverlaysoc_hdmi_in0_chansync_data_out2_de);
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_re = ((~soc_videooverlaysoc_hdmi_in0_chansync_is_control2) | soc_videooverlaysoc_hdmi_in0_chansync_all_control);
assign soc_videooverlaysoc_hdmi_in0_chansync_all_control = ((soc_videooverlaysoc_hdmi_in0_chansync_is_control0 & soc_videooverlaysoc_hdmi_in0_chansync_is_control1) & soc_videooverlaysoc_hdmi_in0_chansync_is_control2);
assign soc_videooverlaysoc_hdmi_in0_chansync_some_control = ((soc_videooverlaysoc_hdmi_in0_chansync_is_control0 | soc_videooverlaysoc_hdmi_in0_chansync_is_control1) | soc_videooverlaysoc_hdmi_in0_chansync_is_control2);
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_adr = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_produce;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_dat_w = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_din;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_we = 1'd1;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_rdport_adr = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_consume;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_dout = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_rdport_dat_r;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_adr = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_produce;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_dat_w = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_din;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_we = 1'd1;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_rdport_adr = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_consume;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_dout = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_rdport_dat_r;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_adr = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_produce;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_dat_w = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_din;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_we = 1'd1;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_rdport_adr = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_consume;
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_dout = soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_rdport_dat_r;
always @(*) begin
	soc_videooverlaysoc_hdmi_in0_decode_terc4_de_o <= 1'd0;
	if (soc_videooverlaysoc_hdmi_in0_decode_terc4_dvimode_bit) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_de_o <= soc_videooverlaysoc_hdmi_in0_decode_terc4_de_r;
	end else begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_de_o <= soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi;
	end
end
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_valid_in = soc_videooverlaysoc_hdmi_in0_decode_terc4_valid_i;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_raw;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_d = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_d;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_c = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_c;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_de = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_de;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_valid_in = soc_videooverlaysoc_hdmi_in0_decode_terc4_valid_i;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_raw;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_d = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_d;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_c = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_c;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_de = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in1_de;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_valid_in = soc_videooverlaysoc_hdmi_in0_decode_terc4_valid_i;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_raw;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_d = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_d;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_c = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_c;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_de = soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in2_de;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_ctl_code = {soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c, soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c};
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_all_vgb = ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb & soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb) & soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb);
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_any_cvalid = ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid | soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid) | soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid);
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_c2c1_dgb = (soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb & soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb);
always @(*) begin
	soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi <= 1'd0;
	vns_clockdomainsrenamer0_next_state0 <= 3'd0;
	soc_videooverlaysoc_hdmi_in0_decode_terc4_encoding_terc4 <= 1'd0;
	soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video <= 1'd0;
	soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data <= 1'd0;
	vns_clockdomainsrenamer0_next_state0 <= vns_clockdomainsrenamer0_state0;
	case (vns_clockdomainsrenamer0_state0)
		1'd1: begin
			if (soc_videooverlaysoc_hdmi_in0_decode_terc4_all_vgb) begin
				vns_clockdomainsrenamer0_next_state0 <= 3'd6;
			end else begin
				if (soc_videooverlaysoc_hdmi_in0_decode_terc4_c2c1_dgb) begin
					vns_clockdomainsrenamer0_next_state0 <= 2'd2;
				end else begin
					if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_ctl_code == 3'd5)) begin
						vns_clockdomainsrenamer0_next_state0 <= 1'd1;
					end else begin
						vns_clockdomainsrenamer0_next_state0 <= 1'd0;
					end
				end
			end
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encoding_terc4 <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi <= 1'd0;
		end
		2'd2: begin
			if (soc_videooverlaysoc_hdmi_in0_decode_terc4_c2c1_dgb) begin
				vns_clockdomainsrenamer0_next_state0 <= 2'd2;
			end else begin
				vns_clockdomainsrenamer0_next_state0 <= 2'd3;
			end
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encoding_terc4 <= 1'd1;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi <= 1'd0;
		end
		2'd3: begin
			if (soc_videooverlaysoc_hdmi_in0_decode_terc4_any_cvalid) begin
				vns_clockdomainsrenamer0_next_state0 <= 1'd0;
			end else begin
				if (soc_videooverlaysoc_hdmi_in0_decode_terc4_all_vgb) begin
					vns_clockdomainsrenamer0_next_state0 <= 3'd6;
				end else begin
					if (soc_videooverlaysoc_hdmi_in0_decode_terc4_c2c1_dgb) begin
						vns_clockdomainsrenamer0_next_state0 <= 3'd4;
					end else begin
						vns_clockdomainsrenamer0_next_state0 <= 2'd3;
					end
				end
			end
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encoding_terc4 <= 1'd1;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data <= 1'd1;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi <= 1'd0;
		end
		3'd4: begin
			if (soc_videooverlaysoc_hdmi_in0_decode_terc4_c2c1_dgb) begin
				vns_clockdomainsrenamer0_next_state0 <= 3'd4;
			end else begin
				vns_clockdomainsrenamer0_next_state0 <= 1'd0;
			end
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encoding_terc4 <= 1'd1;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi <= 1'd0;
		end
		3'd5: begin
			if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_ctl_code == 1'd1)) begin
				vns_clockdomainsrenamer0_next_state0 <= 3'd5;
			end else begin
				if (soc_videooverlaysoc_hdmi_in0_decode_terc4_all_vgb) begin
					vns_clockdomainsrenamer0_next_state0 <= 3'd6;
				end else begin
					vns_clockdomainsrenamer0_next_state0 <= 1'd0;
				end
			end
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encoding_terc4 <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi <= 1'd0;
		end
		3'd6: begin
			if (soc_videooverlaysoc_hdmi_in0_decode_terc4_all_vgb) begin
				vns_clockdomainsrenamer0_next_state0 <= 3'd6;
			end else begin
				vns_clockdomainsrenamer0_next_state0 <= 3'd7;
			end
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encoding_terc4 <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi <= 1'd0;
		end
		3'd7: begin
			if (soc_videooverlaysoc_hdmi_in0_decode_terc4_any_cvalid) begin
				vns_clockdomainsrenamer0_next_state0 <= 1'd0;
			end else begin
				vns_clockdomainsrenamer0_next_state0 <= 3'd7;
			end
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encoding_terc4 <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video <= 1'd1;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi <= 1'd1;
		end
		default: begin
			if (soc_videooverlaysoc_hdmi_in0_decode_terc4_all_vgb) begin
				vns_clockdomainsrenamer0_next_state0 <= 3'd6;
			end else begin
				if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_ctl_code == 3'd5)) begin
					vns_clockdomainsrenamer0_next_state0 <= 1'd1;
				end else begin
					if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_ctl_code == 1'd1)) begin
						vns_clockdomainsrenamer0_next_state0 <= 3'd5;
					end else begin
						vns_clockdomainsrenamer0_next_state0 <= 1'd0;
					end
				end
			end
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encoding_terc4 <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_de_hdmi <= 1'd0;
		end
	endcase
end
assign soc_videooverlaysoc_hdmi_in0_syncpol_de = soc_videooverlaysoc_hdmi_in0_syncpol_de_r;
assign soc_videooverlaysoc_hdmi_in0_syncpol_hsync = soc_videooverlaysoc_hdmi_in0_syncpol_c_out[0];
assign soc_videooverlaysoc_hdmi_in0_syncpol_vsync = soc_videooverlaysoc_hdmi_in0_syncpol_c_out[1];
assign soc_videooverlaysoc_hdmi_in0_syncpol_de_rising = (soc_videooverlaysoc_hdmi_in0_syncpol_de_r & (~soc_videooverlaysoc_hdmi_in0_syncpol_de_int));
assign soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_raw = soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s0;
assign soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_d = soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s1;
assign soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_c = soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s2;
assign soc_videooverlaysoc_hdmi_in0_data0_timingdelay_source_de = soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s3;
assign soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_raw = soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s0;
assign soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_d = soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s1;
assign soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_c = soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s2;
assign soc_videooverlaysoc_hdmi_in0_data1_timingdelay_source_de = soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s3;
assign soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_raw = soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s0;
assign soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_d = soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s1;
assign soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_c = soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s2;
assign soc_videooverlaysoc_hdmi_in0_data2_timingdelay_source_de = soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s3;
assign soc_videooverlaysoc_hdmi_in0_resdetection_pn_de = ((~soc_videooverlaysoc_hdmi_in0_resdetection_de) & soc_videooverlaysoc_hdmi_in0_resdetection_de_r);
assign soc_videooverlaysoc_hdmi_in0_resdetection_p_vsync = (soc_videooverlaysoc_hdmi_in0_resdetection_vsync & (~soc_videooverlaysoc_hdmi_in0_resdetection_vsync_r));
assign soc_videooverlaysoc_hdmi_out0_clk_gen_data1 = (~soc_videooverlaysoc_hdmi_out0_clk_gen_data0);
assign soc_videooverlaysoc_hdmi_out0_phy_sink_ready = 1'd1;
assign soc_videooverlaysoc_hdmi_out0_phy_es0_data0 = soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c0;
assign soc_videooverlaysoc_hdmi_out0_phy_es1_data0 = soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c1;
assign soc_videooverlaysoc_hdmi_out0_phy_es2_data0 = soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c2;
assign soc_videooverlaysoc_hdmi_out0_phy_es0_data1 = soc_videooverlaysoc_hdmi_out0_phy_es0_data0;
assign soc_videooverlaysoc_hdmi_out0_phy_es1_data1 = soc_videooverlaysoc_hdmi_out0_phy_es1_data0;
assign soc_videooverlaysoc_hdmi_out0_phy_es2_data1 = soc_videooverlaysoc_hdmi_out0_phy_es2_data0;
assign hdmi_in1_freq_fmeter_clk = soc_videooverlaysoc_hdmi_in1_freq_clk0;
assign soc_videooverlaysoc_hdmi_in1_freq_period_done = (soc_videooverlaysoc_hdmi_in1_freq_period_counter == 27'd100000000);
assign soc_videooverlaysoc_hdmi_in1_freq_ce = 1'd1;
assign soc_videooverlaysoc_hdmi_in1_freq_sampler_latch = soc_videooverlaysoc_hdmi_in1_freq_period_done;
assign soc_videooverlaysoc_hdmi_in1_freq_sampler_i = soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o;
assign soc_videooverlaysoc_hdmi_in1_freq_status = soc_videooverlaysoc_hdmi_in1_freq_sampler_o;
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_freq_q_next_binary <= 6'd0;
	if (soc_videooverlaysoc_hdmi_in1_freq_ce) begin
		soc_videooverlaysoc_hdmi_in1_freq_q_next_binary <= (soc_videooverlaysoc_hdmi_in1_freq_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_hdmi_in1_freq_q_next_binary <= soc_videooverlaysoc_hdmi_in1_freq_q_binary;
	end
end
assign soc_videooverlaysoc_hdmi_in1_freq_q_next = (soc_videooverlaysoc_hdmi_in1_freq_q_next_binary ^ soc_videooverlaysoc_hdmi_in1_freq_q_next_binary[5:1]);
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb <= 6'd0;
	soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[5] <= soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_i[5];
	soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[4] <= (soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[5] ^ soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_i[4]);
	soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[3] <= (soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[4] ^ soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_i[3]);
	soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[2] <= (soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[3] ^ soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_i[2]);
	soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[1] <= (soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[2] ^ soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_i[1]);
	soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[0] <= (soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb[1] ^ soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_i[0]);
end
assign soc_videooverlaysoc_hdmi_in1_freq_sampler_inc = (soc_videooverlaysoc_hdmi_in1_freq_sampler_i - soc_videooverlaysoc_hdmi_in1_freq_sampler_i_d);
assign soc_videooverlaysoc_hdmi_in1_charsync0_raw_data = soc_videooverlaysoc_hdmi_in1_s7datacapture0_d;
assign soc_videooverlaysoc_hdmi_in1_wer0_data = soc_videooverlaysoc_hdmi_in1_charsync0_data;
assign soc_videooverlaysoc_hdmi_in1_decoding0_valid_i = soc_videooverlaysoc_hdmi_in1_charsync0_synced;
assign soc_videooverlaysoc_hdmi_in1_decoding0_input = soc_videooverlaysoc_hdmi_in1_charsync0_data;
assign soc_videooverlaysoc_hdmi_in1_charsync1_raw_data = soc_videooverlaysoc_hdmi_in1_s7datacapture1_d;
assign soc_videooverlaysoc_hdmi_in1_wer1_data = soc_videooverlaysoc_hdmi_in1_charsync1_data;
assign soc_videooverlaysoc_hdmi_in1_decoding1_valid_i = soc_videooverlaysoc_hdmi_in1_charsync1_synced;
assign soc_videooverlaysoc_hdmi_in1_decoding1_input = soc_videooverlaysoc_hdmi_in1_charsync1_data;
assign soc_videooverlaysoc_hdmi_in1_charsync2_raw_data = soc_videooverlaysoc_hdmi_in1_s7datacapture2_d;
assign soc_videooverlaysoc_hdmi_in1_wer2_data = soc_videooverlaysoc_hdmi_in1_charsync2_data;
assign soc_videooverlaysoc_hdmi_in1_decoding2_valid_i = soc_videooverlaysoc_hdmi_in1_charsync2_synced;
assign soc_videooverlaysoc_hdmi_in1_decoding2_input = soc_videooverlaysoc_hdmi_in1_charsync2_data;
assign soc_videooverlaysoc_hdmi_in1_chansync_valid_i = ((soc_videooverlaysoc_hdmi_in1_decoding0_valid_o & soc_videooverlaysoc_hdmi_in1_decoding1_valid_o) & soc_videooverlaysoc_hdmi_in1_decoding2_valid_o);
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in0_raw = soc_videooverlaysoc_hdmi_in1_decoding0_output_raw;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in0_d = soc_videooverlaysoc_hdmi_in1_decoding0_output_d;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in0_c = soc_videooverlaysoc_hdmi_in1_decoding0_output_c;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in0_de = soc_videooverlaysoc_hdmi_in1_decoding0_output_de;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in1_raw = soc_videooverlaysoc_hdmi_in1_decoding1_output_raw;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in1_d = soc_videooverlaysoc_hdmi_in1_decoding1_output_d;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in1_c = soc_videooverlaysoc_hdmi_in1_decoding1_output_c;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in1_de = soc_videooverlaysoc_hdmi_in1_decoding1_output_de;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in2_raw = soc_videooverlaysoc_hdmi_in1_decoding2_output_raw;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in2_d = soc_videooverlaysoc_hdmi_in1_decoding2_output_d;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in2_c = soc_videooverlaysoc_hdmi_in1_decoding2_output_c;
assign soc_videooverlaysoc_hdmi_in1_chansync_data_in2_de = soc_videooverlaysoc_hdmi_in1_decoding2_output_de;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_valid_i = soc_videooverlaysoc_hdmi_in1_chansync_chan_synced;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_raw = soc_videooverlaysoc_hdmi_in1_chansync_data_out0_raw;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_d = soc_videooverlaysoc_hdmi_in1_chansync_data_out0_d;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_c = soc_videooverlaysoc_hdmi_in1_chansync_data_out0_c;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_de = soc_videooverlaysoc_hdmi_in1_chansync_data_out0_de;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_raw = soc_videooverlaysoc_hdmi_in1_chansync_data_out1_raw;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_d = soc_videooverlaysoc_hdmi_in1_chansync_data_out1_d;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_c = soc_videooverlaysoc_hdmi_in1_chansync_data_out1_c;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_de = soc_videooverlaysoc_hdmi_in1_chansync_data_out1_de;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_raw = soc_videooverlaysoc_hdmi_in1_chansync_data_out2_raw;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_d = soc_videooverlaysoc_hdmi_in1_chansync_data_out2_d;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_c = soc_videooverlaysoc_hdmi_in1_chansync_data_out2_c;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_de = soc_videooverlaysoc_hdmi_in1_chansync_data_out2_de;
assign soc_videooverlaysoc_hdmi_in1_syncpol_de_int = soc_videooverlaysoc_hdmi_in1_decode_terc4_de_o;
assign soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_raw = soc_videooverlaysoc_hdmi_in1_chansync_data_out0_raw;
assign soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_d = soc_videooverlaysoc_hdmi_in1_chansync_data_out0_d;
assign soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_c = soc_videooverlaysoc_hdmi_in1_chansync_data_out0_c;
assign soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_de = soc_videooverlaysoc_hdmi_in1_chansync_data_out0_de;
assign soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_raw = soc_videooverlaysoc_hdmi_in1_chansync_data_out1_raw;
assign soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_d = soc_videooverlaysoc_hdmi_in1_chansync_data_out1_d;
assign soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_c = soc_videooverlaysoc_hdmi_in1_chansync_data_out1_c;
assign soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_de = soc_videooverlaysoc_hdmi_in1_chansync_data_out1_de;
assign soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_raw = soc_videooverlaysoc_hdmi_in1_chansync_data_out2_raw;
assign soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_d = soc_videooverlaysoc_hdmi_in1_chansync_data_out2_d;
assign soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_c = soc_videooverlaysoc_hdmi_in1_chansync_data_out2_c;
assign soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_de = soc_videooverlaysoc_hdmi_in1_chansync_data_out2_de;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_raw = soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_raw;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_d = soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_d;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_c = soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_c;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_de = soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_de;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in1_raw = soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_raw;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in1_d = soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_d;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in1_c = soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_c;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in1_de = soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_de;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in2_raw = soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_raw;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in2_d = soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_d;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in2_c = soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_c;
assign soc_videooverlaysoc_hdmi_in1_syncpol_data_in2_de = soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_de;
assign soc_videooverlaysoc_hdmi_in1_syncpol_valid_i = soc_videooverlaysoc_hdmi_in1_chansync_chan_synced;
assign soc_videooverlaysoc_hdmi_in1_resdetection_valid_i = soc_videooverlaysoc_hdmi_in1_syncpol_valid_o;
assign soc_videooverlaysoc_hdmi_in1_resdetection_de = soc_videooverlaysoc_hdmi_in1_syncpol_de;
assign soc_videooverlaysoc_hdmi_in1_resdetection_vsync = soc_videooverlaysoc_hdmi_in1_syncpol_vsync;
assign soc_videooverlaysoc_hdmi_in1_frame_valid_i = soc_videooverlaysoc_hdmi_in1_syncpol_valid_o;
assign soc_videooverlaysoc_hdmi_in1_frame_de = soc_videooverlaysoc_hdmi_in1_syncpol_de;
assign soc_videooverlaysoc_hdmi_in1_frame_vsync = soc_videooverlaysoc_hdmi_in1_syncpol_vsync;
assign soc_videooverlaysoc_hdmi_in1_frame_r = soc_videooverlaysoc_hdmi_in1_syncpol_r;
assign soc_videooverlaysoc_hdmi_in1_frame_g = soc_videooverlaysoc_hdmi_in1_syncpol_g;
assign soc_videooverlaysoc_hdmi_in1_frame_b = soc_videooverlaysoc_hdmi_in1_syncpol_b;
assign soc_videooverlaysoc_hdmi_in1_dma_frame_valid = soc_videooverlaysoc_hdmi_in1_frame_frame_valid;
assign soc_videooverlaysoc_hdmi_in1_frame_frame_ready = soc_videooverlaysoc_hdmi_in1_dma_frame_ready;
assign soc_videooverlaysoc_hdmi_in1_dma_frame_first = soc_videooverlaysoc_hdmi_in1_frame_frame_first;
assign soc_videooverlaysoc_hdmi_in1_dma_frame_last = soc_videooverlaysoc_hdmi_in1_frame_frame_last;
assign soc_videooverlaysoc_hdmi_in1_dma_frame_payload_sof = soc_videooverlaysoc_hdmi_in1_frame_frame_payload_sof;
assign soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels = soc_videooverlaysoc_hdmi_in1_frame_frame_payload_pixels;
assign soc_videooverlaysoc_hdmi_in1_edid_status = 1'd1;
assign soc_videooverlaysoc_hdmi_in1_edid_sda_o = (~soc_videooverlaysoc_hdmi_in1_edid_sda_drv_reg);
assign soc_videooverlaysoc_hdmi_in1_edid_scl_rising = (soc_videooverlaysoc_hdmi_in1_edid_scl_i & (~soc_videooverlaysoc_hdmi_in1_edid_scl_r));
assign soc_videooverlaysoc_hdmi_in1_edid_sda_rising = (soc_videooverlaysoc_hdmi_in1_edid_sda_i & (~soc_videooverlaysoc_hdmi_in1_edid_sda_r));
assign soc_videooverlaysoc_hdmi_in1_edid_sda_falling = ((~soc_videooverlaysoc_hdmi_in1_edid_sda_i) & soc_videooverlaysoc_hdmi_in1_edid_sda_r);
assign soc_videooverlaysoc_hdmi_in1_edid_start = (soc_videooverlaysoc_hdmi_in1_edid_scl_i & soc_videooverlaysoc_hdmi_in1_edid_sda_falling);
assign soc_videooverlaysoc_hdmi_in1_edid_adr = soc_videooverlaysoc_hdmi_in1_edid_offset_counter;
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_edid_sda_drv <= 1'd0;
	if (soc_videooverlaysoc_hdmi_in1_edid_zero_drv) begin
		soc_videooverlaysoc_hdmi_in1_edid_sda_drv <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_edid_data_drv) begin
			soc_videooverlaysoc_hdmi_in1_edid_sda_drv <= (~soc_videooverlaysoc_hdmi_in1_edid_data_bit);
		end
	end
end
always @(*) begin
	vns_edid1_next_state <= 4'd0;
	soc_videooverlaysoc_hdmi_in1_edid_oc_load <= 1'd0;
	soc_videooverlaysoc_hdmi_in1_edid_oc_inc <= 1'd0;
	soc_videooverlaysoc_hdmi_in1_edid_data_drv_en <= 1'd0;
	soc_videooverlaysoc_hdmi_in1_edid_data_drv_stop <= 1'd0;
	soc_videooverlaysoc_hdmi_in1_edid_update_is_read <= 1'd0;
	soc_videooverlaysoc_hdmi_in1_edid_zero_drv <= 1'd0;
	vns_edid1_next_state <= vns_edid1_state;
	case (vns_edid1_state)
		1'd1: begin
			if ((soc_videooverlaysoc_hdmi_in1_edid_counter == 4'd8)) begin
				if ((soc_videooverlaysoc_hdmi_in1_edid_din[7:1] == 7'd80)) begin
					soc_videooverlaysoc_hdmi_in1_edid_update_is_read <= 1'd1;
					vns_edid1_next_state <= 2'd2;
				end else begin
					vns_edid1_next_state <= 1'd0;
				end
			end
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
		2'd2: begin
			if ((~soc_videooverlaysoc_hdmi_in1_edid_scl_i)) begin
				vns_edid1_next_state <= 2'd3;
			end
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in1_edid_zero_drv <= 1'd1;
			if (soc_videooverlaysoc_hdmi_in1_edid_scl_i) begin
				vns_edid1_next_state <= 3'd4;
			end
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in1_edid_zero_drv <= 1'd1;
			if ((~soc_videooverlaysoc_hdmi_in1_edid_scl_i)) begin
				if (soc_videooverlaysoc_hdmi_in1_edid_is_read) begin
					vns_edid1_next_state <= 4'd9;
				end else begin
					vns_edid1_next_state <= 3'd5;
				end
			end
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
		3'd5: begin
			if ((soc_videooverlaysoc_hdmi_in1_edid_counter == 4'd8)) begin
				soc_videooverlaysoc_hdmi_in1_edid_oc_load <= 1'd1;
				vns_edid1_next_state <= 3'd6;
			end
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
		3'd6: begin
			if ((~soc_videooverlaysoc_hdmi_in1_edid_scl_i)) begin
				vns_edid1_next_state <= 3'd7;
			end
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in1_edid_zero_drv <= 1'd1;
			if (soc_videooverlaysoc_hdmi_in1_edid_scl_i) begin
				vns_edid1_next_state <= 4'd8;
			end
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
		4'd8: begin
			soc_videooverlaysoc_hdmi_in1_edid_zero_drv <= 1'd1;
			if ((~soc_videooverlaysoc_hdmi_in1_edid_scl_i)) begin
				vns_edid1_next_state <= 1'd1;
			end
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
		4'd9: begin
			if ((~soc_videooverlaysoc_hdmi_in1_edid_scl_i)) begin
				if ((soc_videooverlaysoc_hdmi_in1_edid_counter == 4'd8)) begin
					soc_videooverlaysoc_hdmi_in1_edid_data_drv_stop <= 1'd1;
					vns_edid1_next_state <= 4'd10;
				end else begin
					soc_videooverlaysoc_hdmi_in1_edid_data_drv_en <= 1'd1;
				end
			end
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
		4'd10: begin
			if (soc_videooverlaysoc_hdmi_in1_edid_scl_rising) begin
				soc_videooverlaysoc_hdmi_in1_edid_oc_inc <= 1'd1;
				if (soc_videooverlaysoc_hdmi_in1_edid_sda_i) begin
					vns_edid1_next_state <= 1'd0;
				end else begin
					vns_edid1_next_state <= 4'd9;
				end
			end
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
		default: begin
			if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
				vns_edid1_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_hdmi_in1_locked_status = soc_videooverlaysoc_hdmi_in1_locked;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_d = (~soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_q);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_d = soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_q;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i = soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_d = soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_mdata = soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_sdata = soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_d;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_too_late = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_lateness == 8'd255);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_too_early = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_lateness == 1'd0);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_rst = soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_master_inc = soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_master_ce = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_o | soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_o);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_slave_inc = soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_slave_ce = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_o | soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_o);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_r[0]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_r[1]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_r[2]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_r[3]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_r[4]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_reset_lateness = soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_i = soc_videooverlaysoc_hdmi_in1_s7datacapture0_phase_reset_re;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst = (hdmi_in1_pix1p25x_rst | hdmi_in1_pix_rst);
assign hdmi_in1_data0_cap_write_clk = hdmi_in1_pix1p25x_clk;
assign hdmi_in1_data0_cap_read_clk = hdmi_in1_pix_clk;
assign hdmi_in1_data0_cap_write_rst = soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst_write;
assign hdmi_in1_data0_cap_read_rst = soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst_read;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_transition = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_mdata_d != soc_videooverlaysoc_hdmi_in1_s7datacapture0_mdata);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_inc = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_transition & (soc_videooverlaysoc_hdmi_in1_s7datacapture0_mdata == soc_videooverlaysoc_hdmi_in1_s7datacapture0_sdata));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_dec = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_transition & (soc_videooverlaysoc_hdmi_in1_s7datacapture0_mdata != soc_videooverlaysoc_hdmi_in1_s7datacapture0_sdata));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_charsync0_raw = {soc_videooverlaysoc_hdmi_in1_charsync0_raw_data, soc_videooverlaysoc_hdmi_in1_charsync0_raw_data1};
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_wer0_transitions <= 8'd0;
	soc_videooverlaysoc_hdmi_in1_wer0_transitions[0] <= (soc_videooverlaysoc_hdmi_in1_wer0_data_r[0] ^ soc_videooverlaysoc_hdmi_in1_wer0_data_r[1]);
	soc_videooverlaysoc_hdmi_in1_wer0_transitions[1] <= (soc_videooverlaysoc_hdmi_in1_wer0_data_r[1] ^ soc_videooverlaysoc_hdmi_in1_wer0_data_r[2]);
	soc_videooverlaysoc_hdmi_in1_wer0_transitions[2] <= (soc_videooverlaysoc_hdmi_in1_wer0_data_r[2] ^ soc_videooverlaysoc_hdmi_in1_wer0_data_r[3]);
	soc_videooverlaysoc_hdmi_in1_wer0_transitions[3] <= (soc_videooverlaysoc_hdmi_in1_wer0_data_r[3] ^ soc_videooverlaysoc_hdmi_in1_wer0_data_r[4]);
	soc_videooverlaysoc_hdmi_in1_wer0_transitions[4] <= (soc_videooverlaysoc_hdmi_in1_wer0_data_r[4] ^ soc_videooverlaysoc_hdmi_in1_wer0_data_r[5]);
	soc_videooverlaysoc_hdmi_in1_wer0_transitions[5] <= (soc_videooverlaysoc_hdmi_in1_wer0_data_r[5] ^ soc_videooverlaysoc_hdmi_in1_wer0_data_r[6]);
	soc_videooverlaysoc_hdmi_in1_wer0_transitions[6] <= (soc_videooverlaysoc_hdmi_in1_wer0_data_r[6] ^ soc_videooverlaysoc_hdmi_in1_wer0_data_r[7]);
	soc_videooverlaysoc_hdmi_in1_wer0_transitions[7] <= (soc_videooverlaysoc_hdmi_in1_wer0_data_r[7] ^ soc_videooverlaysoc_hdmi_in1_wer0_data_r[8]);
end
assign soc_videooverlaysoc_hdmi_in1_wer0_i = soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_r_updated;
assign soc_videooverlaysoc_hdmi_in1_wer0_o = (soc_videooverlaysoc_hdmi_in1_wer0_toggle_o ^ soc_videooverlaysoc_hdmi_in1_wer0_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_d = soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_q;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_d = (~soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_q);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i = soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_d = soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_mdata = soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_sdata = soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_d;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_too_late = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_lateness == 8'd255);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_too_early = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_lateness == 1'd0);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_rst = soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_master_inc = soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_master_ce = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_o | soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_o);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_slave_inc = soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_slave_ce = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_o | soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_o);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_r[0]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_r[1]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_r[2]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_r[3]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_r[4]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_reset_lateness = soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_i = soc_videooverlaysoc_hdmi_in1_s7datacapture1_phase_reset_re;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst = (hdmi_in1_pix1p25x_rst | hdmi_in1_pix_rst);
assign hdmi_in1_data1_cap_write_clk = hdmi_in1_pix1p25x_clk;
assign hdmi_in1_data1_cap_read_clk = hdmi_in1_pix_clk;
assign hdmi_in1_data1_cap_write_rst = soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst_write;
assign hdmi_in1_data1_cap_read_rst = soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst_read;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_transition = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_mdata_d != soc_videooverlaysoc_hdmi_in1_s7datacapture1_mdata);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_inc = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_transition & (soc_videooverlaysoc_hdmi_in1_s7datacapture1_mdata == soc_videooverlaysoc_hdmi_in1_s7datacapture1_sdata));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_dec = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_transition & (soc_videooverlaysoc_hdmi_in1_s7datacapture1_mdata != soc_videooverlaysoc_hdmi_in1_s7datacapture1_sdata));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_charsync1_raw = {soc_videooverlaysoc_hdmi_in1_charsync1_raw_data, soc_videooverlaysoc_hdmi_in1_charsync1_raw_data1};
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_wer1_transitions <= 8'd0;
	soc_videooverlaysoc_hdmi_in1_wer1_transitions[0] <= (soc_videooverlaysoc_hdmi_in1_wer1_data_r[0] ^ soc_videooverlaysoc_hdmi_in1_wer1_data_r[1]);
	soc_videooverlaysoc_hdmi_in1_wer1_transitions[1] <= (soc_videooverlaysoc_hdmi_in1_wer1_data_r[1] ^ soc_videooverlaysoc_hdmi_in1_wer1_data_r[2]);
	soc_videooverlaysoc_hdmi_in1_wer1_transitions[2] <= (soc_videooverlaysoc_hdmi_in1_wer1_data_r[2] ^ soc_videooverlaysoc_hdmi_in1_wer1_data_r[3]);
	soc_videooverlaysoc_hdmi_in1_wer1_transitions[3] <= (soc_videooverlaysoc_hdmi_in1_wer1_data_r[3] ^ soc_videooverlaysoc_hdmi_in1_wer1_data_r[4]);
	soc_videooverlaysoc_hdmi_in1_wer1_transitions[4] <= (soc_videooverlaysoc_hdmi_in1_wer1_data_r[4] ^ soc_videooverlaysoc_hdmi_in1_wer1_data_r[5]);
	soc_videooverlaysoc_hdmi_in1_wer1_transitions[5] <= (soc_videooverlaysoc_hdmi_in1_wer1_data_r[5] ^ soc_videooverlaysoc_hdmi_in1_wer1_data_r[6]);
	soc_videooverlaysoc_hdmi_in1_wer1_transitions[6] <= (soc_videooverlaysoc_hdmi_in1_wer1_data_r[6] ^ soc_videooverlaysoc_hdmi_in1_wer1_data_r[7]);
	soc_videooverlaysoc_hdmi_in1_wer1_transitions[7] <= (soc_videooverlaysoc_hdmi_in1_wer1_data_r[7] ^ soc_videooverlaysoc_hdmi_in1_wer1_data_r[8]);
end
assign soc_videooverlaysoc_hdmi_in1_wer1_i = soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_r_updated;
assign soc_videooverlaysoc_hdmi_in1_wer1_o = (soc_videooverlaysoc_hdmi_in1_wer1_toggle_o ^ soc_videooverlaysoc_hdmi_in1_wer1_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_d = soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_q;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_d = (~soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_q);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i = soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_d = soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_mdata = soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_d;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_sdata = soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_d;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_too_late = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_lateness == 8'd255);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_too_early = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_lateness == 1'd0);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_rst = soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_master_inc = soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_master_ce = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_o | soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_o);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_slave_inc = soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_slave_ce = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_o | soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_o);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_r[0]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_r[1]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_r[2]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_r[3]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_i = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_re & soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_r[4]);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_reset_lateness = soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_o;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_i = soc_videooverlaysoc_hdmi_in1_s7datacapture2_phase_reset_re;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst = (hdmi_in1_pix1p25x_rst | hdmi_in1_pix_rst);
assign hdmi_in1_data2_cap_write_clk = hdmi_in1_pix1p25x_clk;
assign hdmi_in1_data2_cap_read_clk = hdmi_in1_pix_clk;
assign hdmi_in1_data2_cap_write_rst = soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst_write;
assign hdmi_in1_data2_cap_read_rst = soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst_read;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_transition = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_mdata_d != soc_videooverlaysoc_hdmi_in1_s7datacapture2_mdata);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_inc = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_transition & (soc_videooverlaysoc_hdmi_in1_s7datacapture2_mdata == soc_videooverlaysoc_hdmi_in1_s7datacapture2_sdata));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_dec = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_transition & (soc_videooverlaysoc_hdmi_in1_s7datacapture2_mdata != soc_videooverlaysoc_hdmi_in1_s7datacapture2_sdata));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_o = (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_o ^ soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_charsync2_raw = {soc_videooverlaysoc_hdmi_in1_charsync2_raw_data, soc_videooverlaysoc_hdmi_in1_charsync2_raw_data1};
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_wer2_transitions <= 8'd0;
	soc_videooverlaysoc_hdmi_in1_wer2_transitions[0] <= (soc_videooverlaysoc_hdmi_in1_wer2_data_r[0] ^ soc_videooverlaysoc_hdmi_in1_wer2_data_r[1]);
	soc_videooverlaysoc_hdmi_in1_wer2_transitions[1] <= (soc_videooverlaysoc_hdmi_in1_wer2_data_r[1] ^ soc_videooverlaysoc_hdmi_in1_wer2_data_r[2]);
	soc_videooverlaysoc_hdmi_in1_wer2_transitions[2] <= (soc_videooverlaysoc_hdmi_in1_wer2_data_r[2] ^ soc_videooverlaysoc_hdmi_in1_wer2_data_r[3]);
	soc_videooverlaysoc_hdmi_in1_wer2_transitions[3] <= (soc_videooverlaysoc_hdmi_in1_wer2_data_r[3] ^ soc_videooverlaysoc_hdmi_in1_wer2_data_r[4]);
	soc_videooverlaysoc_hdmi_in1_wer2_transitions[4] <= (soc_videooverlaysoc_hdmi_in1_wer2_data_r[4] ^ soc_videooverlaysoc_hdmi_in1_wer2_data_r[5]);
	soc_videooverlaysoc_hdmi_in1_wer2_transitions[5] <= (soc_videooverlaysoc_hdmi_in1_wer2_data_r[5] ^ soc_videooverlaysoc_hdmi_in1_wer2_data_r[6]);
	soc_videooverlaysoc_hdmi_in1_wer2_transitions[6] <= (soc_videooverlaysoc_hdmi_in1_wer2_data_r[6] ^ soc_videooverlaysoc_hdmi_in1_wer2_data_r[7]);
	soc_videooverlaysoc_hdmi_in1_wer2_transitions[7] <= (soc_videooverlaysoc_hdmi_in1_wer2_data_r[7] ^ soc_videooverlaysoc_hdmi_in1_wer2_data_r[8]);
end
assign soc_videooverlaysoc_hdmi_in1_wer2_i = soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_r_updated;
assign soc_videooverlaysoc_hdmi_in1_wer2_o = (soc_videooverlaysoc_hdmi_in1_wer2_toggle_o ^ soc_videooverlaysoc_hdmi_in1_wer2_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_din = {soc_videooverlaysoc_hdmi_in1_chansync_data_in0_de, soc_videooverlaysoc_hdmi_in1_chansync_data_in0_c, soc_videooverlaysoc_hdmi_in1_chansync_data_in0_d, soc_videooverlaysoc_hdmi_in1_chansync_data_in0_raw};
assign {soc_videooverlaysoc_hdmi_in1_chansync_data_out0_de, soc_videooverlaysoc_hdmi_in1_chansync_data_out0_c, soc_videooverlaysoc_hdmi_in1_chansync_data_out0_d, soc_videooverlaysoc_hdmi_in1_chansync_data_out0_raw} = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_dout;
assign soc_videooverlaysoc_hdmi_in1_chansync_is_control0 = (~soc_videooverlaysoc_hdmi_in1_chansync_data_out0_de);
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_re = ((~soc_videooverlaysoc_hdmi_in1_chansync_is_control0) | soc_videooverlaysoc_hdmi_in1_chansync_all_control);
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_din = {soc_videooverlaysoc_hdmi_in1_chansync_data_in1_de, soc_videooverlaysoc_hdmi_in1_chansync_data_in1_c, soc_videooverlaysoc_hdmi_in1_chansync_data_in1_d, soc_videooverlaysoc_hdmi_in1_chansync_data_in1_raw};
assign {soc_videooverlaysoc_hdmi_in1_chansync_data_out1_de, soc_videooverlaysoc_hdmi_in1_chansync_data_out1_c, soc_videooverlaysoc_hdmi_in1_chansync_data_out1_d, soc_videooverlaysoc_hdmi_in1_chansync_data_out1_raw} = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_dout;
assign soc_videooverlaysoc_hdmi_in1_chansync_is_control1 = (~soc_videooverlaysoc_hdmi_in1_chansync_data_out1_de);
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_re = ((~soc_videooverlaysoc_hdmi_in1_chansync_is_control1) | soc_videooverlaysoc_hdmi_in1_chansync_all_control);
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_din = {soc_videooverlaysoc_hdmi_in1_chansync_data_in2_de, soc_videooverlaysoc_hdmi_in1_chansync_data_in2_c, soc_videooverlaysoc_hdmi_in1_chansync_data_in2_d, soc_videooverlaysoc_hdmi_in1_chansync_data_in2_raw};
assign {soc_videooverlaysoc_hdmi_in1_chansync_data_out2_de, soc_videooverlaysoc_hdmi_in1_chansync_data_out2_c, soc_videooverlaysoc_hdmi_in1_chansync_data_out2_d, soc_videooverlaysoc_hdmi_in1_chansync_data_out2_raw} = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_dout;
assign soc_videooverlaysoc_hdmi_in1_chansync_is_control2 = (~soc_videooverlaysoc_hdmi_in1_chansync_data_out2_de);
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_re = ((~soc_videooverlaysoc_hdmi_in1_chansync_is_control2) | soc_videooverlaysoc_hdmi_in1_chansync_all_control);
assign soc_videooverlaysoc_hdmi_in1_chansync_all_control = ((soc_videooverlaysoc_hdmi_in1_chansync_is_control0 & soc_videooverlaysoc_hdmi_in1_chansync_is_control1) & soc_videooverlaysoc_hdmi_in1_chansync_is_control2);
assign soc_videooverlaysoc_hdmi_in1_chansync_some_control = ((soc_videooverlaysoc_hdmi_in1_chansync_is_control0 | soc_videooverlaysoc_hdmi_in1_chansync_is_control1) | soc_videooverlaysoc_hdmi_in1_chansync_is_control2);
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_adr = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_produce;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_dat_w = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_din;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_we = 1'd1;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_rdport_adr = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_consume;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_dout = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_rdport_dat_r;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_adr = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_produce;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_dat_w = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_din;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_we = 1'd1;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_rdport_adr = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_consume;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_dout = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_rdport_dat_r;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_adr = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_produce;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_dat_w = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_din;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_we = 1'd1;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_rdport_adr = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_consume;
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_dout = soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_rdport_dat_r;
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_decode_terc4_de_o <= 1'd0;
	if (soc_videooverlaysoc_hdmi_in1_decode_terc4_dvimode_bit) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_de_o <= soc_videooverlaysoc_hdmi_in1_decode_terc4_de_r;
	end else begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_de_o <= soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi;
	end
end
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_valid_in = soc_videooverlaysoc_hdmi_in1_decode_terc4_valid_i;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_raw;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_d = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_d;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_c = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_c;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_de = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_de;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_valid_in = soc_videooverlaysoc_hdmi_in1_decode_terc4_valid_i;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_raw;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_d = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_d;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_c = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_c;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_de = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in1_de;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_valid_in = soc_videooverlaysoc_hdmi_in1_decode_terc4_valid_i;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_raw;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_d = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_d;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_c = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_c;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_de = soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in2_de;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_ctl_code = {soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c, soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c};
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_all_vgb = ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb & soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb) & soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb);
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_any_cvalid = ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid | soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid) | soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid);
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_c2c1_dgb = (soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb & soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb);
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi <= 1'd0;
	soc_videooverlaysoc_hdmi_in1_decode_terc4_encoding_terc4 <= 1'd0;
	vns_clockdomainsrenamer1_next_state0 <= 3'd0;
	soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_video <= 1'd0;
	soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_data <= 1'd0;
	vns_clockdomainsrenamer1_next_state0 <= vns_clockdomainsrenamer1_state0;
	case (vns_clockdomainsrenamer1_state0)
		1'd1: begin
			if (soc_videooverlaysoc_hdmi_in1_decode_terc4_all_vgb) begin
				vns_clockdomainsrenamer1_next_state0 <= 3'd6;
			end else begin
				if (soc_videooverlaysoc_hdmi_in1_decode_terc4_c2c1_dgb) begin
					vns_clockdomainsrenamer1_next_state0 <= 2'd2;
				end else begin
					if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_ctl_code == 3'd5)) begin
						vns_clockdomainsrenamer1_next_state0 <= 1'd1;
					end else begin
						vns_clockdomainsrenamer1_next_state0 <= 1'd0;
					end
				end
			end
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encoding_terc4 <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi <= 1'd0;
		end
		2'd2: begin
			if (soc_videooverlaysoc_hdmi_in1_decode_terc4_c2c1_dgb) begin
				vns_clockdomainsrenamer1_next_state0 <= 2'd2;
			end else begin
				vns_clockdomainsrenamer1_next_state0 <= 2'd3;
			end
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encoding_terc4 <= 1'd1;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi <= 1'd0;
		end
		2'd3: begin
			if (soc_videooverlaysoc_hdmi_in1_decode_terc4_any_cvalid) begin
				vns_clockdomainsrenamer1_next_state0 <= 1'd0;
			end else begin
				if (soc_videooverlaysoc_hdmi_in1_decode_terc4_all_vgb) begin
					vns_clockdomainsrenamer1_next_state0 <= 3'd6;
				end else begin
					if (soc_videooverlaysoc_hdmi_in1_decode_terc4_c2c1_dgb) begin
						vns_clockdomainsrenamer1_next_state0 <= 3'd4;
					end else begin
						vns_clockdomainsrenamer1_next_state0 <= 2'd3;
					end
				end
			end
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encoding_terc4 <= 1'd1;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_data <= 1'd1;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi <= 1'd0;
		end
		3'd4: begin
			if (soc_videooverlaysoc_hdmi_in1_decode_terc4_c2c1_dgb) begin
				vns_clockdomainsrenamer1_next_state0 <= 3'd4;
			end else begin
				vns_clockdomainsrenamer1_next_state0 <= 1'd0;
			end
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encoding_terc4 <= 1'd1;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi <= 1'd0;
		end
		3'd5: begin
			if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_ctl_code == 1'd1)) begin
				vns_clockdomainsrenamer1_next_state0 <= 3'd5;
			end else begin
				if (soc_videooverlaysoc_hdmi_in1_decode_terc4_all_vgb) begin
					vns_clockdomainsrenamer1_next_state0 <= 3'd6;
				end else begin
					vns_clockdomainsrenamer1_next_state0 <= 1'd0;
				end
			end
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encoding_terc4 <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi <= 1'd0;
		end
		3'd6: begin
			if (soc_videooverlaysoc_hdmi_in1_decode_terc4_all_vgb) begin
				vns_clockdomainsrenamer1_next_state0 <= 3'd6;
			end else begin
				vns_clockdomainsrenamer1_next_state0 <= 3'd7;
			end
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encoding_terc4 <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi <= 1'd0;
		end
		3'd7: begin
			if (soc_videooverlaysoc_hdmi_in1_decode_terc4_any_cvalid) begin
				vns_clockdomainsrenamer1_next_state0 <= 1'd0;
			end else begin
				vns_clockdomainsrenamer1_next_state0 <= 3'd7;
			end
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encoding_terc4 <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_video <= 1'd1;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi <= 1'd1;
		end
		default: begin
			if (soc_videooverlaysoc_hdmi_in1_decode_terc4_all_vgb) begin
				vns_clockdomainsrenamer1_next_state0 <= 3'd6;
			end else begin
				if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_ctl_code == 3'd5)) begin
					vns_clockdomainsrenamer1_next_state0 <= 1'd1;
				end else begin
					if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_ctl_code == 1'd1)) begin
						vns_clockdomainsrenamer1_next_state0 <= 3'd5;
					end else begin
						vns_clockdomainsrenamer1_next_state0 <= 1'd0;
					end
				end
			end
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encoding_terc4 <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_data <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_encrypting_video <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_de_hdmi <= 1'd0;
		end
	endcase
end
assign soc_videooverlaysoc_hdmi_in1_syncpol_de = soc_videooverlaysoc_hdmi_in1_syncpol_de_r;
assign soc_videooverlaysoc_hdmi_in1_syncpol_hsync = soc_videooverlaysoc_hdmi_in1_syncpol_c_out[0];
assign soc_videooverlaysoc_hdmi_in1_syncpol_vsync = soc_videooverlaysoc_hdmi_in1_syncpol_c_out[1];
assign soc_videooverlaysoc_hdmi_in1_syncpol_de_rising = (soc_videooverlaysoc_hdmi_in1_syncpol_de_r & (~soc_videooverlaysoc_hdmi_in1_syncpol_de_int));
assign soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_raw = soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s0;
assign soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_d = soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s1;
assign soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_c = soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s2;
assign soc_videooverlaysoc_hdmi_in1_data0_timingdelay_source_de = soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s3;
assign soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_raw = soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s0;
assign soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_d = soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s1;
assign soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_c = soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s2;
assign soc_videooverlaysoc_hdmi_in1_data1_timingdelay_source_de = soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s3;
assign soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_raw = soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s0;
assign soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_d = soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s1;
assign soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_c = soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s2;
assign soc_videooverlaysoc_hdmi_in1_data2_timingdelay_source_de = soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s3;
assign soc_videooverlaysoc_hdmi_in1_resdetection_pn_de = ((~soc_videooverlaysoc_hdmi_in1_resdetection_de) & soc_videooverlaysoc_hdmi_in1_resdetection_de_r);
assign soc_videooverlaysoc_hdmi_in1_resdetection_p_vsync = (soc_videooverlaysoc_hdmi_in1_resdetection_vsync & (~soc_videooverlaysoc_hdmi_in1_resdetection_vsync_r));
assign soc_videooverlaysoc_hdmi_in1_frame_new_frame = (soc_videooverlaysoc_hdmi_in1_frame_vsync & (~soc_videooverlaysoc_hdmi_in1_frame_vsync_r));
assign soc_videooverlaysoc_hdmi_in1_frame_encoded_pixel = {soc_videooverlaysoc_hdmi_in1_frame_dummy8, soc_videooverlaysoc_hdmi_in1_frame_r, soc_videooverlaysoc_hdmi_in1_frame_g, soc_videooverlaysoc_hdmi_in1_frame_b};
assign soc_videooverlaysoc_hdmi_in1_frame_sink_payload_pixels = soc_videooverlaysoc_hdmi_in1_frame_cur_word;
assign soc_videooverlaysoc_hdmi_in1_frame_sink_valid = soc_videooverlaysoc_hdmi_in1_frame_cur_word_valid;
assign soc_videooverlaysoc_hdmi_in1_frame_frame_valid = soc_videooverlaysoc_hdmi_in1_frame_source_valid;
assign soc_videooverlaysoc_hdmi_in1_frame_source_ready = soc_videooverlaysoc_hdmi_in1_frame_frame_ready;
assign soc_videooverlaysoc_hdmi_in1_frame_frame_first = soc_videooverlaysoc_hdmi_in1_frame_source_first;
assign soc_videooverlaysoc_hdmi_in1_frame_frame_last = soc_videooverlaysoc_hdmi_in1_frame_source_last;
assign soc_videooverlaysoc_hdmi_in1_frame_frame_payload_sof = soc_videooverlaysoc_hdmi_in1_frame_source_payload_sof;
assign soc_videooverlaysoc_hdmi_in1_frame_frame_payload_pixels = soc_videooverlaysoc_hdmi_in1_frame_source_payload_pixels;
assign soc_videooverlaysoc_hdmi_in1_frame_busy = 1'd0;
assign soc_videooverlaysoc_hdmi_in1_frame_pix_overflow_reset = soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_o;
assign soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_i = soc_videooverlaysoc_hdmi_in1_frame_pix_overflow_reset;
assign soc_videooverlaysoc_hdmi_in1_frame_overflow_w = (soc_videooverlaysoc_hdmi_in1_frame_sys_overflow & (~soc_videooverlaysoc_hdmi_in1_frame_overflow_mask));
assign soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_i = soc_videooverlaysoc_hdmi_in1_frame_overflow_re;
assign soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_din = {soc_videooverlaysoc_hdmi_in1_frame_fifo_in_last, soc_videooverlaysoc_hdmi_in1_frame_fifo_in_first, soc_videooverlaysoc_hdmi_in1_frame_fifo_in_payload_pixels, soc_videooverlaysoc_hdmi_in1_frame_fifo_in_payload_sof};
assign {soc_videooverlaysoc_hdmi_in1_frame_fifo_out_last, soc_videooverlaysoc_hdmi_in1_frame_fifo_out_first, soc_videooverlaysoc_hdmi_in1_frame_fifo_out_payload_pixels, soc_videooverlaysoc_hdmi_in1_frame_fifo_out_payload_sof} = soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_dout;
assign soc_videooverlaysoc_hdmi_in1_frame_sink_ready = soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_writable;
assign soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_we = soc_videooverlaysoc_hdmi_in1_frame_sink_valid;
assign soc_videooverlaysoc_hdmi_in1_frame_fifo_in_first = soc_videooverlaysoc_hdmi_in1_frame_sink_first;
assign soc_videooverlaysoc_hdmi_in1_frame_fifo_in_last = soc_videooverlaysoc_hdmi_in1_frame_sink_last;
assign soc_videooverlaysoc_hdmi_in1_frame_fifo_in_payload_sof = soc_videooverlaysoc_hdmi_in1_frame_sink_payload_sof;
assign soc_videooverlaysoc_hdmi_in1_frame_fifo_in_payload_pixels = soc_videooverlaysoc_hdmi_in1_frame_sink_payload_pixels;
assign soc_videooverlaysoc_hdmi_in1_frame_source_valid = soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_readable;
assign soc_videooverlaysoc_hdmi_in1_frame_source_first = soc_videooverlaysoc_hdmi_in1_frame_fifo_out_first;
assign soc_videooverlaysoc_hdmi_in1_frame_source_last = soc_videooverlaysoc_hdmi_in1_frame_fifo_out_last;
assign soc_videooverlaysoc_hdmi_in1_frame_source_payload_sof = soc_videooverlaysoc_hdmi_in1_frame_fifo_out_payload_sof;
assign soc_videooverlaysoc_hdmi_in1_frame_source_payload_pixels = soc_videooverlaysoc_hdmi_in1_frame_fifo_out_payload_pixels;
assign soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_re = soc_videooverlaysoc_hdmi_in1_frame_source_ready;
assign soc_videooverlaysoc_hdmi_in1_frame_graycounter0_ce = (soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_writable & soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_we);
assign soc_videooverlaysoc_hdmi_in1_frame_graycounter1_ce = (soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_readable & soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_re);
assign soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_writable = (((soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q[10] == soc_videooverlaysoc_hdmi_in1_frame_consume_wdomain[10]) | (soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q[9] == soc_videooverlaysoc_hdmi_in1_frame_consume_wdomain[9])) | (soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q[8:0] != soc_videooverlaysoc_hdmi_in1_frame_consume_wdomain[8:0]));
assign soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_readable = (soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q != soc_videooverlaysoc_hdmi_in1_frame_produce_rdomain);
assign soc_videooverlaysoc_hdmi_in1_frame_wrport_adr = soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_binary[9:0];
assign soc_videooverlaysoc_hdmi_in1_frame_wrport_dat_w = soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_din;
assign soc_videooverlaysoc_hdmi_in1_frame_wrport_we = soc_videooverlaysoc_hdmi_in1_frame_graycounter0_ce;
assign soc_videooverlaysoc_hdmi_in1_frame_rdport_adr = soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next_binary[9:0];
assign soc_videooverlaysoc_hdmi_in1_frame_asyncfifo_dout = soc_videooverlaysoc_hdmi_in1_frame_rdport_dat_r;
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_next_binary <= 11'd0;
	if (soc_videooverlaysoc_hdmi_in1_frame_graycounter0_ce) begin
		soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_next_binary <= (soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_next_binary <= soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_binary;
	end
end
assign soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_next = (soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_next_binary ^ soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_next_binary[10:1]);
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next_binary <= 11'd0;
	if (soc_videooverlaysoc_hdmi_in1_frame_graycounter1_ce) begin
		soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next_binary <= (soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next_binary <= soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_binary;
	end
end
assign soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next = (soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next_binary ^ soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next_binary[10:1]);
assign soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_o = (soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_o ^ soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_o = (soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_o ^ soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_o_r);
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_reached = soc_videooverlaysoc_hdmi_in1_dma_current_address;
assign soc_videooverlaysoc_hdmi_in1_dma_last_word = (soc_videooverlaysoc_hdmi_in1_dma_mwords_remaining == 1'd1);
assign soc_videooverlaysoc_hdmi_in1_dma_memory_word = {soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels, soc_videooverlaysoc_hdmi_in1_dma_frame_payload_pixels};
assign soc_videooverlaysoc_hdmi_in1_dma_sink_sink_payload_address = soc_videooverlaysoc_hdmi_in1_dma_current_address;
assign soc_videooverlaysoc_hdmi_in1_dma_sink_sink_payload_data = soc_videooverlaysoc_hdmi_in1_dma_memory_word;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_change_slot = ((~soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_valid) | soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_done);
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_address = vns_comb_rhs_array_muxed36;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_valid = vns_comb_rhs_array_muxed37;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_reached = soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_reached;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_reached = soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_reached;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_done = (soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_done & (soc_videooverlaysoc_hdmi_in1_dma_slot_array_current_slot == 1'd0));
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_done = (soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_done & (soc_videooverlaysoc_hdmi_in1_dma_slot_array_current_slot == 1'd1));
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_clear <= 1'd0;
	if ((soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_re & soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_r[0])) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_clear <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_status_w <= 2'd0;
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_status_w[0] <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status;
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_status_w[1] <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status;
end
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_clear <= 1'd0;
	if ((soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_re & soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_r[1])) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_clear <= 1'd1;
	end
end
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_w <= 2'd0;
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_w[0] <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_pending;
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_w[1] <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_pending;
end
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_irq = ((soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_w[0] & soc_videooverlaysoc_hdmi_in1_dma_slot_array_storage[0]) | (soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_w[1] & soc_videooverlaysoc_hdmi_in1_dma_slot_array_storage[1]));
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_trigger;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_pending = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_trigger;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_trigger;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_pending = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_trigger;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_valid = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_storage[0];
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_dat_w = 2'd2;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_we = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_done;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_dat_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_reached;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_we = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_done;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_trigger = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_storage[1];
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_valid = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_storage[0];
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_dat_w = 2'd2;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_we = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_done;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_dat_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_reached;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_we = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_done;
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_trigger = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_storage[1];
assign soc_videooverlaysoc_litedramcrossbar_cmd_payload_we = 1'd1;
assign soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr = soc_videooverlaysoc_hdmi_in1_dma_sink_sink_payload_address;
assign soc_videooverlaysoc_litedramcrossbar_cmd_valid = (soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_ready & soc_videooverlaysoc_hdmi_in1_dma_sink_sink_valid);
assign soc_videooverlaysoc_hdmi_in1_dma_sink_sink_ready = (soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_ready & soc_videooverlaysoc_litedramcrossbar_cmd_ready);
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_valid = (soc_videooverlaysoc_hdmi_in1_dma_sink_sink_valid & soc_videooverlaysoc_litedramcrossbar_cmd_ready);
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_payload_data = soc_videooverlaysoc_hdmi_in1_dma_sink_sink_payload_data;
assign soc_videooverlaysoc_litedramcrossbar_wdata_payload_we = 32'd4294967295;
assign soc_videooverlaysoc_litedramcrossbar_wdata_valid = soc_videooverlaysoc_hdmi_in1_dma_fifo_source_valid;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_source_ready = soc_videooverlaysoc_litedramcrossbar_wdata_ready;
assign soc_videooverlaysoc_litedramcrossbar_wdata_payload_data = soc_videooverlaysoc_hdmi_in1_dma_fifo_source_payload_data;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_din = {soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_in_last, soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_in_first, soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_in_payload_data};
assign {soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_out_last, soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_out_first, soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_out_payload_data} = soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_dout;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_ready = soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_writable;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_we = soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_valid;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_in_first = soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_first;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_in_last = soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_last;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_in_payload_data = soc_videooverlaysoc_hdmi_in1_dma_fifo_sink_payload_data;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_source_valid = soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_readable;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_source_first = soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_out_first;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_source_last = soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_out_last;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_source_payload_data = soc_videooverlaysoc_hdmi_in1_dma_fifo_fifo_out_payload_data;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_re = soc_videooverlaysoc_hdmi_in1_dma_fifo_source_ready;
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_adr <= 4'd0;
	if (soc_videooverlaysoc_hdmi_in1_dma_fifo_replace) begin
		soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_adr <= (soc_videooverlaysoc_hdmi_in1_dma_fifo_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_adr <= soc_videooverlaysoc_hdmi_in1_dma_fifo_produce;
	end
end
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_dat_w = soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_din;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_we = (soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_we & (soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_writable | soc_videooverlaysoc_hdmi_in1_dma_fifo_replace));
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_do_read = (soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_readable & soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_re);
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_rdport_adr = soc_videooverlaysoc_hdmi_in1_dma_fifo_consume;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_dout = soc_videooverlaysoc_hdmi_in1_dma_fifo_rdport_dat_r;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_writable = (soc_videooverlaysoc_hdmi_in1_dma_fifo_level != 5'd16);
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_readable = (soc_videooverlaysoc_hdmi_in1_dma_fifo_level != 1'd0);
always @(*) begin
	soc_videooverlaysoc_hdmi_in1_dma_count_word <= 1'd0;
	soc_videooverlaysoc_hdmi_in1_dma_sink_sink_valid <= 1'd0;
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_done <= 1'd0;
	soc_videooverlaysoc_hdmi_in1_dma_frame_ready <= 1'd0;
	vns_dma_next_state <= 2'd0;
	soc_videooverlaysoc_hdmi_in1_dma_reset_words <= 1'd0;
	vns_dma_next_state <= vns_dma_state;
	case (vns_dma_state)
		1'd1: begin
			soc_videooverlaysoc_hdmi_in1_dma_frame_ready <= soc_videooverlaysoc_hdmi_in1_dma_sink_sink_ready;
			if (soc_videooverlaysoc_hdmi_in1_dma_frame_valid) begin
				soc_videooverlaysoc_hdmi_in1_dma_sink_sink_valid <= 1'd1;
				if (soc_videooverlaysoc_hdmi_in1_dma_sink_sink_ready) begin
					soc_videooverlaysoc_hdmi_in1_dma_count_word <= 1'd1;
					if (soc_videooverlaysoc_hdmi_in1_dma_last_word) begin
						vns_dma_next_state <= 2'd2;
					end
				end
			end
		end
		2'd2: begin
			if ((~soc_videooverlaysoc_litedramcrossbar_wdata_valid)) begin
				soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_done <= 1'd1;
				vns_dma_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_hdmi_in1_dma_reset_words <= 1'd1;
			soc_videooverlaysoc_hdmi_in1_dma_frame_ready <= ((~soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_valid) | (~soc_videooverlaysoc_hdmi_in1_dma_frame_payload_sof));
			if (((soc_videooverlaysoc_hdmi_in1_dma_slot_array_address_valid & soc_videooverlaysoc_hdmi_in1_dma_frame_payload_sof) & soc_videooverlaysoc_hdmi_in1_dma_frame_valid)) begin
				vns_dma_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_valid = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_valid;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_valid = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_valid;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_ready = soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_ready;
assign soc_videooverlaysoc_hdmi_core_out0_source_source_valid = (soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_valid & ((~soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_de) | soc_videooverlaysoc_hdmi_core_out0_dmareader_source_valid));
always @(*) begin
	soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_ready <= 1'd0;
	soc_videooverlaysoc_hdmi_core_out0_dmareader_source_ready <= 1'd0;
	if ((~soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_valid)) begin
		soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_ready <= 1'd1;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_source_ready <= 1'd1;
	end else begin
		if ((soc_videooverlaysoc_hdmi_core_out0_source_source_valid & soc_videooverlaysoc_hdmi_core_out0_source_source_ready)) begin
			soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_ready <= 1'd1;
			soc_videooverlaysoc_hdmi_core_out0_dmareader_source_ready <= (soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_de | 1'd0);
		end
	end
end
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_hres = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hres;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_hsync_start = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hsync_start;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_hsync_end = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hsync_end;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_hscan = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hscan;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_vres = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vres;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_vsync_start = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vsync_start;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_vsync_end = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vsync_end;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_sink_payload_vscan = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vscan;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_payload_base = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_base;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_payload_length = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_length;
assign soc_videooverlaysoc_hdmi_core_out0_source_source_param_de = soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_de;
assign soc_videooverlaysoc_hdmi_core_out0_source_source_param_hsync = soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_hsync;
assign soc_videooverlaysoc_hdmi_core_out0_source_source_param_vsync = soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_vsync;
assign soc_videooverlaysoc_hdmi_core_out0_source_source_payload_data = soc_videooverlaysoc_hdmi_core_out0_dmareader_source_payload_data;
assign soc_videooverlaysoc_hdmi_core_out0_i = soc_videooverlaysoc_hdmi_core_out0_underflow_update_underflow_update_re;
assign soc_videooverlaysoc_hdmi_core_out0_underflow_update = soc_videooverlaysoc_hdmi_core_out0_o;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hres = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hsync_start = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hsync_end = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hscan = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vres = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vsync_start = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vsync_end = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vscan = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_base = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_length = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_valid = soc_videooverlaysoc_hdmi_core_out0_initiator_enable_storage;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_valid = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_valid;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_ready = soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_ready;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_first = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_first;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_last = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_last;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hres = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hres;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hsync_start = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hsync_start;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hsync_end = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hsync_end;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_hscan = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hscan;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vres = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vres;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vsync_start = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vsync_start;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vsync_end = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vsync_end;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_vscan = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vscan;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_base = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_base;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_source_source_payload_length = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_length;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_din = {soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_last, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_first, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_length, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_base, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vscan, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vsync_end, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vsync_start, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vres, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hscan, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hsync_end, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hsync_start, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hres};
assign {soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_last, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_first, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_length, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_base, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vscan, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vsync_end, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vsync_start, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vres, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hscan, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hsync_end, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hsync_start, soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hres} = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_dout;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_ready = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_writable;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_we = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_valid;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_first = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_first;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_last = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_last;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hres = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hres;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hsync_start = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hsync_start;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hsync_end = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hsync_end;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_hscan = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_hscan;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vres = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vres;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vsync_start = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vsync_start;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vsync_end = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vsync_end;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_vscan = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_vscan;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_base = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_base;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_in_payload_length = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_sink_payload_length;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_valid = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_readable;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_first = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_first;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_last = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_last;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hres = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hres;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hsync_start = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hsync_start;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hsync_end = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hsync_end;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_hscan = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_hscan;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vres = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vres;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vsync_start = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vsync_start;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vsync_end = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vsync_end;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_vscan = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_vscan;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_base = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_base;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_payload_length = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_fifo_out_payload_length;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_re = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_source_ready;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_ce = (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_writable & soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_we);
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_ce = (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_readable & soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_re);
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_writable = ((soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q[1] == soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_consume_wdomain[1]) | (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q[0] == soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_consume_wdomain[0]));
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_readable = (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q != soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_produce_rdomain);
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_adr = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_binary[0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_dat_w = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_din;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_we = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_ce;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_rdport_adr = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next_binary[0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_asyncfifo_dout = soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_rdport_dat_r;
always @(*) begin
	soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_next_binary <= 2'd0;
	if (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_ce) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_next_binary <= (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_next_binary <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_binary;
	end
end
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_next = (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_next_binary ^ soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_next_binary[1]);
always @(*) begin
	soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next_binary <= 2'd0;
	if (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_ce) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next_binary <= (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next_binary <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_binary;
	end
end
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next = (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next_binary ^ soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next_binary[1]);
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_valid = soc_videooverlaysoc_hdmi_in0_timing_valid;
assign soc_videooverlaysoc_hdmi_in0_timing_ready = soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_ready;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_first = soc_videooverlaysoc_hdmi_in0_timing_first;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_last = soc_videooverlaysoc_hdmi_in0_timing_last;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_hsync = soc_videooverlaysoc_hdmi_in0_timing_payload_hsync;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_vsync = soc_videooverlaysoc_hdmi_in0_timing_payload_vsync;
assign soc_videooverlaysoc_hdmi_core_out0_timinggenerator_source_payload_de = soc_videooverlaysoc_hdmi_in0_timing_payload_de;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_base = soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_payload_base[31:2];
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_length = soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_payload_length[31:2];
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_sink_payload_address = (soc_videooverlaysoc_hdmi_core_out0_dmareader_base + soc_videooverlaysoc_hdmi_core_out0_dmareader_offset);
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_source_valid = soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_valid;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_ready = soc_videooverlaysoc_hdmi_core_out0_dmareader_source_ready;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_source_first = soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_first;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_source_last = soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_last;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_source_payload_data = soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_payload_data;
assign soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_payload_we = 1'd0;
assign soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_payload_addr = soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_sink_payload_address;
assign soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_valid = (soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_sink_valid & soc_videooverlaysoc_hdmi_core_out0_dmareader_request_enable);
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_sink_ready = (soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_ready & soc_videooverlaysoc_hdmi_core_out0_dmareader_request_enable);
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_request_issued = (soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_valid & soc_videooverlaysoc_out_dram_port_litedramnativeport1_cmd_ready);
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_request_enable = (soc_videooverlaysoc_hdmi_core_out0_dmareader_rsv_level != 11'd1024);
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_valid = soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_valid;
assign soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_ready = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_ready;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_first = soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_first;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_last = soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_last;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_payload_data = soc_videooverlaysoc_out_dram_port_litedramnativeport1_rdata_payload_data;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_valid = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_valid;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_ready = soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_ready;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_first = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_first;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_last = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_last;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_payload_data = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_payload_data;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_data_dequeued = (soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_valid & soc_videooverlaysoc_hdmi_core_out0_dmareader_source_source_ready);
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_din = {soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_in_last, soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_in_first, soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_in_payload_data};
assign {soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_out_last, soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_out_first, soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_out_payload_data} = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_dout;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_ready = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_writable;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_we = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_valid;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_in_first = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_first;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_in_last = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_last;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_in_payload_data = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_sink_payload_data;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_valid = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_readable;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_first = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_out_first;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_last = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_out_last;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_payload_data = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_fifo_out_payload_data;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_re = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_source_ready;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_re = (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_readable & ((~soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_readable) | soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_re));
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level1 = (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level0 + soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_readable);
always @(*) begin
	soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_adr <= 10'd0;
	if (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_replace) begin
		soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_adr <= (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_adr <= soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_produce;
	end
end
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_dat_w = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_din;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_we = (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_we & (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_writable | soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_replace));
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_do_read = (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_readable & soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_re);
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_rdport_adr = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_consume;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_dout = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_rdport_dat_r;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_rdport_re = soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_do_read;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_writable = (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level0 != 11'd1024);
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_readable = (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level0 != 1'd0);
always @(*) begin
	vns_videooutcore_next_state <= 2'd0;
	soc_videooverlaysoc_hdmi_core_out0_dmareader_offset_next_value <= 27'd0;
	soc_videooverlaysoc_hdmi_core_out0_dmareader_offset_next_value_ce <= 1'd0;
	soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_ready <= 1'd0;
	soc_videooverlaysoc_out_dram_port_litedramnativeport1_flush <= 1'd0;
	soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_sink_valid <= 1'd0;
	vns_videooutcore_next_state <= vns_videooutcore_state;
	case (vns_videooutcore_state)
		1'd1: begin
			soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_sink_valid <= 1'd1;
			if (soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_sink_ready) begin
				soc_videooverlaysoc_hdmi_core_out0_dmareader_offset_next_value <= (soc_videooverlaysoc_hdmi_core_out0_dmareader_offset + 1'd1);
				soc_videooverlaysoc_hdmi_core_out0_dmareader_offset_next_value_ce <= 1'd1;
				if ((soc_videooverlaysoc_hdmi_core_out0_dmareader_offset == (soc_videooverlaysoc_hdmi_core_out0_dmareader_length - 1'd1))) begin
					soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_ready <= 1'd1;
					vns_videooutcore_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			if (soc_videooverlaysoc_hdmi_core_out0_dmareader_sof) begin
				vns_videooutcore_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_hdmi_core_out0_dmareader_offset_next_value <= soc_videooverlaysoc_hdmi_core_out0_dmareader_storage;
			soc_videooverlaysoc_hdmi_core_out0_dmareader_offset_next_value_ce <= 1'd1;
			if (soc_videooverlaysoc_hdmi_core_out0_dmareader_sink_valid) begin
				vns_videooutcore_next_state <= 1'd1;
			end else begin
				soc_videooverlaysoc_out_dram_port_litedramnativeport1_flush <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_hdmi_core_out0_o = (soc_videooverlaysoc_hdmi_core_out0_toggle_o ^ soc_videooverlaysoc_hdmi_core_out0_toggle_o_r);
assign soc_videooverlaysoc_timing_rgb_delay_source_payload_r = soc_videooverlaysoc_timing_rgb_delay_next_s3;
assign soc_videooverlaysoc_timing_rgb_delay_source_payload_g = soc_videooverlaysoc_timing_rgb_delay_next_s7;
assign soc_videooverlaysoc_timing_rgb_delay_source_payload_b = soc_videooverlaysoc_timing_rgb_delay_next_s11;
assign soc_videooverlaysoc_i2c_snoop_status = soc_videooverlaysoc_i2c_snoop_reg_dout;
assign soc_videooverlaysoc_encoder0_q_m8_n = ((soc_videooverlaysoc_encoder0_n1d > 3'd4) | ((soc_videooverlaysoc_encoder0_n1d == 3'd4) & (~soc_videooverlaysoc_encoder0_d1[0])));
assign soc_videooverlaysoc_encoder1_q_m8_n = ((soc_videooverlaysoc_encoder1_n1d > 3'd4) | ((soc_videooverlaysoc_encoder1_n1d == 3'd4) & (~soc_videooverlaysoc_encoder1_d1[0])));
assign soc_videooverlaysoc_encoder2_q_m8_n = ((soc_videooverlaysoc_encoder2_n1d > 3'd4) | ((soc_videooverlaysoc_encoder2_n1d == 3'd4) & (~soc_videooverlaysoc_encoder2_d1[0])));
assign soc_videooverlaysoc_rect_on1 = (((((soc_videooverlaysoc_hcounter > soc_videooverlaysoc_hrect_start_storage) & (soc_videooverlaysoc_hcounter < soc_videooverlaysoc_hrect_end_storage)) & (soc_videooverlaysoc_vcounter > soc_videooverlaysoc_vrect_start_storage)) & (soc_videooverlaysoc_vcounter < soc_videooverlaysoc_vrect_end_storage)) == 1'd1);
assign eth_rx_clk = eth_clk;
assign eth_tx_clk = eth_clk;
assign soc_videooverlaysoc_phy_reset0 = (soc_videooverlaysoc_phy_reset_storage | soc_videooverlaysoc_phy_reset1);
assign rmii_eth_rst_n = (~soc_videooverlaysoc_phy_reset0);
assign soc_videooverlaysoc_phy_counter_done = (soc_videooverlaysoc_phy_counter == 9'd256);
assign soc_videooverlaysoc_phy_counter_ce = (~soc_videooverlaysoc_phy_counter_done);
assign soc_videooverlaysoc_phy_reset1 = (~soc_videooverlaysoc_phy_counter_done);
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_valid = soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_valid;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_payload_data = soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_payload_data;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_ready = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_ready;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_ready = 1'd1;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_valid = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_valid;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_first = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_first;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_last = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_last;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_ready = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_ready;
always @(*) begin
	soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_payload_data <= 8'd0;
	soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_payload_data[1:0] <= soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_payload_data[1:0];
	soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_payload_data[3:2] <= soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_payload_data[3:2];
	soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_payload_data[5:4] <= soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_payload_data[5:4];
	soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_payload_data[7:6] <= soc_videooverlaysoc_phy_liteethphyrmiitx_converter_sink_payload_data[7:6];
end
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_valid = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_valid;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_first = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_first;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_last = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_last;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_ready = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_ready;
assign {soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_payload_data} = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_payload_data;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_valid = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_valid;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_ready = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_ready;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_first = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_first;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_last = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_last;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_source_payload_data = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_payload_data;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_first = (soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_mux == 1'd0);
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_last = (soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_mux == 2'd3);
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_valid = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_valid;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_first = (soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_first & soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_first);
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_last = (soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_last & soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_last);
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_ready = (soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_last & soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_ready);
always @(*) begin
	soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_payload_data <= 2'd0;
	case (soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_mux)
		1'd0: begin
			soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_payload_data <= soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_payload_data[1:0];
		end
		1'd1: begin
			soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_payload_data <= soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_payload_data[3:2];
		end
		2'd2: begin
			soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_payload_data <= soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_payload_data[5:4];
		end
		default: begin
			soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_payload_data <= soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_sink_payload_data[7:6];
		end
	endcase
end
assign soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_payload_valid_token_count = soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_last;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_valid = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_valid;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_ready = soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_ready;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_first = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_first;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_last = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_last;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_payload_data = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_payload_data;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_valid = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_valid0;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_first = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_first;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_last = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_last;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_ready = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_ready;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_payload_data = {soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_payload_data};
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_valid = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_valid;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_first = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_first;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_last = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_last;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_ready = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_ready;
always @(*) begin
	soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_payload_data <= 8'd0;
	soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_payload_data[1:0] <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_payload_data[1:0];
	soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_payload_data[3:2] <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_payload_data[3:2];
	soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_payload_data[5:4] <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_payload_data[5:4];
	soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_payload_data[7:6] <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_payload_data[7:6];
end
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_valid = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_valid;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_ready = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_ready;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_first = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_first;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_last = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_last;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_source_source_payload_data = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_data;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_ready = ((~soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_strobe_all) | soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_ready);
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_valid = soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_strobe_all;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_load_part = (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_valid & soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_ready);
always @(*) begin
	soc_videooverlaysoc_phy_liteethphyrmiirx_converter_reset <= 1'd0;
	soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_valid1 <= 1'd0;
	vns_clockdomainsrenamer0_next_state1 <= 1'd0;
	soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_data <= 2'd0;
	soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_last <= 1'd0;
	vns_clockdomainsrenamer0_next_state1 <= vns_clockdomainsrenamer0_state1;
	case (vns_clockdomainsrenamer0_state1)
		1'd1: begin
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_valid1 <= 1'd1;
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_data <= soc_videooverlaysoc_phy_liteethphyrmiirx_rx_data;
			if ((~(soc_videooverlaysoc_phy_liteethphyrmiirx_crs_dv | soc_videooverlaysoc_phy_liteethphyrmiirx_crs_dv_d))) begin
				soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_last <= 1'd1;
				vns_clockdomainsrenamer0_next_state1 <= 1'd0;
			end
		end
		default: begin
			if ((soc_videooverlaysoc_phy_liteethphyrmiirx_crs_dv & (soc_videooverlaysoc_phy_liteethphyrmiirx_rx_data != 1'd0))) begin
				soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_valid1 <= 1'd1;
				soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_data <= soc_videooverlaysoc_phy_liteethphyrmiirx_rx_data;
				vns_clockdomainsrenamer0_next_state1 <= 1'd1;
			end else begin
				soc_videooverlaysoc_phy_liteethphyrmiirx_converter_reset <= 1'd1;
			end
		end
	endcase
end
assign rmii_eth_mdc = soc_videooverlaysoc_phy_storage[0];
assign soc_videooverlaysoc_phy_data_oe = soc_videooverlaysoc_phy_storage[1];
assign soc_videooverlaysoc_phy_data_w = soc_videooverlaysoc_phy_storage[2];
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_valid = soc_videooverlaysoc_core_mac_crossbar_source_valid;
assign soc_videooverlaysoc_core_mac_crossbar_source_ready = soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_ready;
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_first = soc_videooverlaysoc_core_mac_crossbar_source_first;
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_last = soc_videooverlaysoc_core_mac_crossbar_source_last;
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_ethernet_type = soc_videooverlaysoc_core_mac_crossbar_source_payload_ethernet_type;
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_sender_mac = soc_videooverlaysoc_core_mac_crossbar_source_payload_sender_mac;
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_target_mac = soc_videooverlaysoc_core_mac_crossbar_source_payload_target_mac;
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_data = soc_videooverlaysoc_core_mac_crossbar_source_payload_data;
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_last_be = soc_videooverlaysoc_core_mac_crossbar_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_error = soc_videooverlaysoc_core_mac_crossbar_source_payload_error;
assign soc_videooverlaysoc_core_mac_tx_cdc_sink_valid = soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_valid;
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_ready = soc_videooverlaysoc_core_mac_tx_cdc_sink_ready;
assign soc_videooverlaysoc_core_mac_tx_cdc_sink_first = soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_first;
assign soc_videooverlaysoc_core_mac_tx_cdc_sink_last = soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_last;
assign soc_videooverlaysoc_core_mac_tx_cdc_sink_payload_data = soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_data;
assign soc_videooverlaysoc_core_mac_tx_cdc_sink_payload_last_be = soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_tx_cdc_sink_payload_error = soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_error;
assign soc_videooverlaysoc_core_mac_depacketizer_sink_valid = soc_videooverlaysoc_core_mac_rx_cdc_source_valid;
assign soc_videooverlaysoc_core_mac_rx_cdc_source_ready = soc_videooverlaysoc_core_mac_depacketizer_sink_ready;
assign soc_videooverlaysoc_core_mac_depacketizer_sink_first = soc_videooverlaysoc_core_mac_rx_cdc_source_first;
assign soc_videooverlaysoc_core_mac_depacketizer_sink_last = soc_videooverlaysoc_core_mac_rx_cdc_source_last;
assign soc_videooverlaysoc_core_mac_depacketizer_sink_payload_data = soc_videooverlaysoc_core_mac_rx_cdc_source_payload_data;
assign soc_videooverlaysoc_core_mac_depacketizer_sink_payload_last_be = soc_videooverlaysoc_core_mac_rx_cdc_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_depacketizer_sink_payload_error = soc_videooverlaysoc_core_mac_rx_cdc_source_payload_error;
assign soc_videooverlaysoc_core_mac_crossbar_sink_valid = soc_videooverlaysoc_core_mac_depacketizer_source_valid;
assign soc_videooverlaysoc_core_mac_depacketizer_source_ready = soc_videooverlaysoc_core_mac_crossbar_sink_ready;
assign soc_videooverlaysoc_core_mac_crossbar_sink_first = soc_videooverlaysoc_core_mac_depacketizer_source_first;
assign soc_videooverlaysoc_core_mac_crossbar_sink_last = soc_videooverlaysoc_core_mac_depacketizer_source_last;
assign soc_videooverlaysoc_core_mac_crossbar_sink_payload_ethernet_type = soc_videooverlaysoc_core_mac_depacketizer_source_payload_ethernet_type;
assign soc_videooverlaysoc_core_mac_crossbar_sink_payload_sender_mac = soc_videooverlaysoc_core_mac_depacketizer_source_payload_sender_mac;
assign soc_videooverlaysoc_core_mac_crossbar_sink_payload_target_mac = soc_videooverlaysoc_core_mac_depacketizer_source_payload_target_mac;
assign soc_videooverlaysoc_core_mac_crossbar_sink_payload_data = soc_videooverlaysoc_core_mac_depacketizer_source_payload_data;
assign soc_videooverlaysoc_core_mac_crossbar_sink_payload_last_be = soc_videooverlaysoc_core_mac_depacketizer_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_crossbar_sink_payload_error = soc_videooverlaysoc_core_mac_depacketizer_source_payload_error;
assign soc_videooverlaysoc_core_mac_ps_preamble_error_i = soc_videooverlaysoc_core_mac_preamble_checker_error;
assign soc_videooverlaysoc_core_mac_ps_crc_error_i = soc_videooverlaysoc_core_mac_crc32_checker_error;
always @(*) begin
	soc_videooverlaysoc_core_mac_tx_gap_inserter_source_valid <= 1'd0;
	soc_videooverlaysoc_core_mac_tx_gap_inserter_source_first <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmacgap_next_state <= 1'd0;
	soc_videooverlaysoc_core_mac_tx_gap_inserter_source_last <= 1'd0;
	soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_last_be <= 1'd0;
	soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_mac_tx_gap_inserter_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_mac_tx_gap_inserter_counter_ce <= 1'd0;
	soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_ready <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmacgap_next_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacgap_state;
	case (vns_clockdomainsrenamer1_liteethmac_liteethmacgap_state)
		1'd1: begin
			soc_videooverlaysoc_core_mac_tx_gap_inserter_counter_ce <= 1'd1;
			if ((soc_videooverlaysoc_core_mac_tx_gap_inserter_counter == 4'd11)) begin
				vns_clockdomainsrenamer1_liteethmac_liteethmacgap_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_mac_tx_gap_inserter_counter_reset <= 1'd1;
			soc_videooverlaysoc_core_mac_tx_gap_inserter_source_valid <= soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_valid;
			soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_ready <= soc_videooverlaysoc_core_mac_tx_gap_inserter_source_ready;
			soc_videooverlaysoc_core_mac_tx_gap_inserter_source_first <= soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_first;
			soc_videooverlaysoc_core_mac_tx_gap_inserter_source_last <= soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_last;
			soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_payload_data;
			soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_last_be <= soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_payload_last_be;
			soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_error <= soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_payload_error;
			if (((soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_valid & soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_last) & soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_ready)) begin
				vns_clockdomainsrenamer1_liteethmac_liteethmacgap_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_last_be = soc_videooverlaysoc_core_mac_preamble_inserter_sink_payload_last_be;
always @(*) begin
	soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_inserter_clr_cnt <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_inserter_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_inserter_inc_cnt <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_next_state <= 2'd0;
	soc_videooverlaysoc_core_mac_preamble_inserter_source_valid <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_inserter_source_first <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_inserter_source_last <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_preamble_inserter_sink_payload_data;
	vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_next_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_state;
	case (vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_state)
		1'd1: begin
			soc_videooverlaysoc_core_mac_preamble_inserter_source_valid <= 1'd1;
			case (soc_videooverlaysoc_core_mac_preamble_inserter_cnt)
				1'd0: begin
					soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_preamble_inserter_preamble[7:0];
				end
				1'd1: begin
					soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_preamble_inserter_preamble[15:8];
				end
				2'd2: begin
					soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_preamble_inserter_preamble[23:16];
				end
				2'd3: begin
					soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_preamble_inserter_preamble[31:24];
				end
				3'd4: begin
					soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_preamble_inserter_preamble[39:32];
				end
				3'd5: begin
					soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_preamble_inserter_preamble[47:40];
				end
				3'd6: begin
					soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_preamble_inserter_preamble[55:48];
				end
				default: begin
					soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_preamble_inserter_preamble[63:56];
				end
			endcase
			if ((soc_videooverlaysoc_core_mac_preamble_inserter_cnt == 3'd7)) begin
				if (soc_videooverlaysoc_core_mac_preamble_inserter_source_ready) begin
					vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_next_state <= 2'd2;
				end
			end else begin
				soc_videooverlaysoc_core_mac_preamble_inserter_inc_cnt <= soc_videooverlaysoc_core_mac_preamble_inserter_source_ready;
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_mac_preamble_inserter_source_valid <= soc_videooverlaysoc_core_mac_preamble_inserter_sink_valid;
			soc_videooverlaysoc_core_mac_preamble_inserter_sink_ready <= soc_videooverlaysoc_core_mac_preamble_inserter_source_ready;
			soc_videooverlaysoc_core_mac_preamble_inserter_source_first <= soc_videooverlaysoc_core_mac_preamble_inserter_sink_first;
			soc_videooverlaysoc_core_mac_preamble_inserter_source_last <= soc_videooverlaysoc_core_mac_preamble_inserter_sink_last;
			soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_error <= soc_videooverlaysoc_core_mac_preamble_inserter_sink_payload_error;
			if (((soc_videooverlaysoc_core_mac_preamble_inserter_sink_valid & soc_videooverlaysoc_core_mac_preamble_inserter_sink_last) & soc_videooverlaysoc_core_mac_preamble_inserter_source_ready)) begin
				vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_mac_preamble_inserter_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_mac_preamble_inserter_clr_cnt <= 1'd1;
			if (soc_videooverlaysoc_core_mac_preamble_inserter_sink_valid) begin
				soc_videooverlaysoc_core_mac_preamble_inserter_sink_ready <= 1'd0;
				vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_mac_preamble_checker_source_payload_data = soc_videooverlaysoc_core_mac_preamble_checker_sink_payload_data;
assign soc_videooverlaysoc_core_mac_preamble_checker_source_payload_last_be = soc_videooverlaysoc_core_mac_preamble_checker_sink_payload_last_be;
always @(*) begin
	soc_videooverlaysoc_core_mac_preamble_checker_error <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_checker_source_valid <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_checker_source_last <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_checker_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_checker_source_first <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_next_state <= 1'd0;
	soc_videooverlaysoc_core_mac_preamble_checker_source_payload_error <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_next_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_state;
	case (vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_state)
		1'd1: begin
			soc_videooverlaysoc_core_mac_preamble_checker_source_valid <= soc_videooverlaysoc_core_mac_preamble_checker_sink_valid;
			soc_videooverlaysoc_core_mac_preamble_checker_sink_ready <= soc_videooverlaysoc_core_mac_preamble_checker_source_ready;
			soc_videooverlaysoc_core_mac_preamble_checker_source_first <= soc_videooverlaysoc_core_mac_preamble_checker_sink_first;
			soc_videooverlaysoc_core_mac_preamble_checker_source_last <= soc_videooverlaysoc_core_mac_preamble_checker_sink_last;
			soc_videooverlaysoc_core_mac_preamble_checker_source_payload_error <= soc_videooverlaysoc_core_mac_preamble_checker_sink_payload_error;
			if (((soc_videooverlaysoc_core_mac_preamble_checker_source_valid & soc_videooverlaysoc_core_mac_preamble_checker_source_last) & soc_videooverlaysoc_core_mac_preamble_checker_source_ready)) begin
				vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_mac_preamble_checker_sink_ready <= 1'd1;
			if (((soc_videooverlaysoc_core_mac_preamble_checker_sink_valid & (~soc_videooverlaysoc_core_mac_preamble_checker_sink_last)) & (soc_videooverlaysoc_core_mac_preamble_checker_sink_payload_data == 8'd213))) begin
				vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_next_state <= 1'd1;
			end
			if ((soc_videooverlaysoc_core_mac_preamble_checker_sink_valid & soc_videooverlaysoc_core_mac_preamble_checker_sink_last)) begin
				soc_videooverlaysoc_core_mac_preamble_checker_error <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_mac_crc32_inserter_cnt_done = (soc_videooverlaysoc_core_mac_crc32_inserter_cnt == 1'd0);
assign soc_videooverlaysoc_core_mac_crc32_inserter_data1 = soc_videooverlaysoc_core_mac_crc32_inserter_data0;
assign soc_videooverlaysoc_core_mac_crc32_inserter_last = soc_videooverlaysoc_core_mac_crc32_inserter_reg;
assign soc_videooverlaysoc_core_mac_crc32_inserter_value = (~{soc_videooverlaysoc_core_mac_crc32_inserter_reg[0], soc_videooverlaysoc_core_mac_crc32_inserter_reg[1], soc_videooverlaysoc_core_mac_crc32_inserter_reg[2], soc_videooverlaysoc_core_mac_crc32_inserter_reg[3], soc_videooverlaysoc_core_mac_crc32_inserter_reg[4], soc_videooverlaysoc_core_mac_crc32_inserter_reg[5], soc_videooverlaysoc_core_mac_crc32_inserter_reg[6], soc_videooverlaysoc_core_mac_crc32_inserter_reg[7], soc_videooverlaysoc_core_mac_crc32_inserter_reg[8], soc_videooverlaysoc_core_mac_crc32_inserter_reg[9], soc_videooverlaysoc_core_mac_crc32_inserter_reg[10], soc_videooverlaysoc_core_mac_crc32_inserter_reg[11], soc_videooverlaysoc_core_mac_crc32_inserter_reg[12], soc_videooverlaysoc_core_mac_crc32_inserter_reg[13], soc_videooverlaysoc_core_mac_crc32_inserter_reg[14], soc_videooverlaysoc_core_mac_crc32_inserter_reg[15], soc_videooverlaysoc_core_mac_crc32_inserter_reg[16], soc_videooverlaysoc_core_mac_crc32_inserter_reg[17], soc_videooverlaysoc_core_mac_crc32_inserter_reg[18], soc_videooverlaysoc_core_mac_crc32_inserter_reg[19], soc_videooverlaysoc_core_mac_crc32_inserter_reg[20], soc_videooverlaysoc_core_mac_crc32_inserter_reg[21], soc_videooverlaysoc_core_mac_crc32_inserter_reg[22], soc_videooverlaysoc_core_mac_crc32_inserter_reg[23], soc_videooverlaysoc_core_mac_crc32_inserter_reg[24], soc_videooverlaysoc_core_mac_crc32_inserter_reg[25], soc_videooverlaysoc_core_mac_crc32_inserter_reg[26], soc_videooverlaysoc_core_mac_crc32_inserter_reg[27], soc_videooverlaysoc_core_mac_crc32_inserter_reg[28], soc_videooverlaysoc_core_mac_crc32_inserter_reg[29], soc_videooverlaysoc_core_mac_crc32_inserter_reg[30], soc_videooverlaysoc_core_mac_crc32_inserter_reg[31]});
assign soc_videooverlaysoc_core_mac_crc32_inserter_error = (soc_videooverlaysoc_core_mac_crc32_inserter_next != 32'd3338984827);
always @(*) begin
	soc_videooverlaysoc_core_mac_crc32_inserter_next <= 32'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_next[0] <= (((soc_videooverlaysoc_core_mac_crc32_inserter_last[24] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[1] <= (((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[25] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[2] <= (((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[26] ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[3] <= (((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[27] ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[4] <= (((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[28] ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[5] <= (((((((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[29] ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[6] <= (((((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[30] ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[7] <= (((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[31] ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[8] <= ((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[0] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[9] <= ((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[1] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[10] <= ((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[2] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[11] <= ((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[3] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[12] <= ((((((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[4] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[13] <= ((((((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[5] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[14] <= ((((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[6] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[15] <= ((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[7] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[16] <= ((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[8] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[17] <= ((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[9] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[18] <= ((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[10] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[19] <= ((((soc_videooverlaysoc_core_mac_crc32_inserter_last[11] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[20] <= ((soc_videooverlaysoc_core_mac_crc32_inserter_last[12] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[21] <= ((soc_videooverlaysoc_core_mac_crc32_inserter_last[13] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[22] <= ((soc_videooverlaysoc_core_mac_crc32_inserter_last[14] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[23] <= ((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[15] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[24] <= ((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[16] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[25] <= ((((soc_videooverlaysoc_core_mac_crc32_inserter_last[17] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[26] <= ((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[18] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[27] <= ((((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[19] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[28] <= ((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[20] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[5]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[29] <= ((((((soc_videooverlaysoc_core_mac_crc32_inserter_last[21] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[4]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[30] <= ((((soc_videooverlaysoc_core_mac_crc32_inserter_last[22] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[3]);
	soc_videooverlaysoc_core_mac_crc32_inserter_next[31] <= ((soc_videooverlaysoc_core_mac_crc32_inserter_last[23] ^ soc_videooverlaysoc_core_mac_crc32_inserter_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_inserter_data1[2]);
end
always @(*) begin
	soc_videooverlaysoc_core_mac_crc32_inserter_source_last <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_last_be <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_data0 <= 8'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_is_ongoing0 <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_is_ongoing1 <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_ce <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_reset <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_source_valid <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_next_state <= 2'd0;
	soc_videooverlaysoc_core_mac_crc32_inserter_source_first <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_next_state <= vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_state;
	case (vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_state)
		1'd1: begin
			soc_videooverlaysoc_core_mac_crc32_inserter_ce <= (soc_videooverlaysoc_core_mac_crc32_inserter_sink_valid & soc_videooverlaysoc_core_mac_crc32_inserter_source_ready);
			soc_videooverlaysoc_core_mac_crc32_inserter_data0 <= soc_videooverlaysoc_core_mac_crc32_inserter_sink_payload_data;
			soc_videooverlaysoc_core_mac_crc32_inserter_source_valid <= soc_videooverlaysoc_core_mac_crc32_inserter_sink_valid;
			soc_videooverlaysoc_core_mac_crc32_inserter_sink_ready <= soc_videooverlaysoc_core_mac_crc32_inserter_source_ready;
			soc_videooverlaysoc_core_mac_crc32_inserter_source_first <= soc_videooverlaysoc_core_mac_crc32_inserter_sink_first;
			soc_videooverlaysoc_core_mac_crc32_inserter_source_last <= soc_videooverlaysoc_core_mac_crc32_inserter_sink_last;
			soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_crc32_inserter_sink_payload_data;
			soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_last_be <= soc_videooverlaysoc_core_mac_crc32_inserter_sink_payload_last_be;
			soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_error <= soc_videooverlaysoc_core_mac_crc32_inserter_sink_payload_error;
			soc_videooverlaysoc_core_mac_crc32_inserter_source_last <= 1'd0;
			if (((soc_videooverlaysoc_core_mac_crc32_inserter_sink_valid & soc_videooverlaysoc_core_mac_crc32_inserter_sink_last) & soc_videooverlaysoc_core_mac_crc32_inserter_source_ready)) begin
				vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_mac_crc32_inserter_source_valid <= 1'd1;
			case (soc_videooverlaysoc_core_mac_crc32_inserter_cnt)
				1'd0: begin
					soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_crc32_inserter_value[31:24];
				end
				1'd1: begin
					soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_crc32_inserter_value[23:16];
				end
				2'd2: begin
					soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_crc32_inserter_value[15:8];
				end
				default: begin
					soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_crc32_inserter_value[7:0];
				end
			endcase
			if (soc_videooverlaysoc_core_mac_crc32_inserter_cnt_done) begin
				soc_videooverlaysoc_core_mac_crc32_inserter_source_last <= 1'd1;
				if (soc_videooverlaysoc_core_mac_crc32_inserter_source_ready) begin
					vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_next_state <= 1'd0;
				end
			end
			soc_videooverlaysoc_core_mac_crc32_inserter_is_ongoing1 <= 1'd1;
		end
		default: begin
			soc_videooverlaysoc_core_mac_crc32_inserter_reset <= 1'd1;
			soc_videooverlaysoc_core_mac_crc32_inserter_sink_ready <= 1'd1;
			if (soc_videooverlaysoc_core_mac_crc32_inserter_sink_valid) begin
				soc_videooverlaysoc_core_mac_crc32_inserter_sink_ready <= 1'd0;
				vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_next_state <= 1'd1;
			end
			soc_videooverlaysoc_core_mac_crc32_inserter_is_ongoing0 <= 1'd1;
		end
	endcase
end
assign soc_videooverlaysoc_core_mac_crc32_checker_fifo_full = (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_level == 3'd4);
assign soc_videooverlaysoc_core_mac_crc32_checker_fifo_in = (soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_valid & ((~soc_videooverlaysoc_core_mac_crc32_checker_fifo_full) | soc_videooverlaysoc_core_mac_crc32_checker_fifo_out));
assign soc_videooverlaysoc_core_mac_crc32_checker_fifo_out = (soc_videooverlaysoc_core_mac_crc32_checker_source_source_valid & soc_videooverlaysoc_core_mac_crc32_checker_source_source_ready);
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_first = soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_first;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_last = soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_last;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_payload_data = soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_data;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_payload_last_be = soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_last_be;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_payload_error = soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_error;
always @(*) begin
	soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_valid <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_valid <= soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_valid;
	soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_valid <= soc_videooverlaysoc_core_mac_crc32_checker_fifo_in;
end
always @(*) begin
	soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_ready <= soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_ready;
	soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_ready <= soc_videooverlaysoc_core_mac_crc32_checker_fifo_in;
end
assign soc_videooverlaysoc_core_mac_crc32_checker_source_source_valid = (soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_valid & soc_videooverlaysoc_core_mac_crc32_checker_fifo_full);
assign soc_videooverlaysoc_core_mac_crc32_checker_source_source_last = soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_last;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_ready = soc_videooverlaysoc_core_mac_crc32_checker_fifo_out;
assign soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_data = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_payload_data;
assign soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_last_be = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_payload_last_be;
always @(*) begin
	soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_error <= soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_payload_error;
	soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_error <= (soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_error | soc_videooverlaysoc_core_mac_crc32_checker_crc_error);
end
assign soc_videooverlaysoc_core_mac_crc32_checker_error = ((soc_videooverlaysoc_core_mac_crc32_checker_source_source_valid & soc_videooverlaysoc_core_mac_crc32_checker_source_source_last) & soc_videooverlaysoc_core_mac_crc32_checker_crc_error);
assign soc_videooverlaysoc_core_mac_crc32_checker_crc_data0 = soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_data;
assign soc_videooverlaysoc_core_mac_crc32_checker_crc_data1 = soc_videooverlaysoc_core_mac_crc32_checker_crc_data0;
assign soc_videooverlaysoc_core_mac_crc32_checker_crc_last = soc_videooverlaysoc_core_mac_crc32_checker_crc_reg;
assign soc_videooverlaysoc_core_mac_crc32_checker_crc_value = (~{soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[0], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[1], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[2], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[3], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[4], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[5], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[6], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[7], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[8], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[9], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[10], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[11], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[12], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[13], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[14], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[15], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[16], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[17], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[18], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[19], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[20], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[21], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[22], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[23], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[24], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[25], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[26], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[27], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[28], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[29], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[30], soc_videooverlaysoc_core_mac_crc32_checker_crc_reg[31]});
assign soc_videooverlaysoc_core_mac_crc32_checker_crc_error = (soc_videooverlaysoc_core_mac_crc32_checker_crc_next != 32'd3338984827);
always @(*) begin
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next <= 32'd0;
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[0] <= (((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[1] <= (((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[2] <= (((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[3] <= (((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[4] <= (((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[5] <= (((((((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[6] <= (((((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[7] <= (((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[8] <= ((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[0] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[9] <= ((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[1] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[10] <= ((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[2] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[11] <= ((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[3] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[12] <= ((((((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[4] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[13] <= ((((((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[5] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[14] <= ((((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[6] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[15] <= ((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[7] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[16] <= ((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[8] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[17] <= ((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[9] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[18] <= ((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[10] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[19] <= ((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[11] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[20] <= ((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[12] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[21] <= ((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[13] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[22] <= ((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[14] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[23] <= ((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[15] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[24] <= ((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[16] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[25] <= ((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[17] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[26] <= ((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[18] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[24]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[7]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[27] <= ((((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[19] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[25]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[6]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[28] <= ((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[20] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[26]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[5]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[29] <= ((((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[21] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[30]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[1]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[27]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[4]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[30] <= ((((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[22] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[31]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[0]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[28]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[3]);
	soc_videooverlaysoc_core_mac_crc32_checker_crc_next[31] <= ((soc_videooverlaysoc_core_mac_crc32_checker_crc_last[23] ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_last[29]) ^ soc_videooverlaysoc_core_mac_crc32_checker_crc_data1[2]);
end
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_din = {soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_last, soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_first, soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_payload_error, soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_payload_last_be, soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_payload_data};
assign {soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_last, soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_first, soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_payload_error, soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_payload_last_be, soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_payload_data} = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_dout;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_ready = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_writable;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_we = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_valid;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_first = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_first;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_last = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_last;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_payload_data = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_payload_data;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_payload_last_be = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_payload_last_be;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_in_payload_error = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_sink_payload_error;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_valid = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_readable;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_first = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_first;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_last = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_last;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_payload_data = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_payload_data;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_payload_last_be = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_payload_last_be;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_payload_error = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_fifo_out_payload_error;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_re = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_source_ready;
always @(*) begin
	soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_adr <= 3'd0;
	if (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_replace) begin
		soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_adr <= (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_adr <= soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_produce;
	end
end
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_dat_w = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_din;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_we = (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_we & (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_writable | soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_replace));
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_do_read = (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_readable & soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_re);
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_rdport_adr = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_consume;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_dout = soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_rdport_dat_r;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_writable = (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_level != 3'd5);
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_readable = (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_level != 1'd0);
always @(*) begin
	vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_next_state <= 2'd0;
	soc_videooverlaysoc_core_mac_crc32_checker_crc_reset <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_checker_fifo_reset <= 1'd0;
	soc_videooverlaysoc_core_mac_crc32_checker_crc_ce <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_next_state <= vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_state;
	case (vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_state)
		1'd1: begin
			if ((soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_valid & soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_ready)) begin
				soc_videooverlaysoc_core_mac_crc32_checker_crc_ce <= 1'd1;
				vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if ((soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_valid & soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_ready)) begin
				soc_videooverlaysoc_core_mac_crc32_checker_crc_ce <= 1'd1;
				if (soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_last) begin
					vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_core_mac_crc32_checker_crc_reset <= 1'd1;
			soc_videooverlaysoc_core_mac_crc32_checker_fifo_reset <= 1'd1;
			vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_next_state <= 1'd1;
		end
	endcase
end
assign soc_videooverlaysoc_core_mac_ps_preamble_error_o = (soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_o ^ soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_o_r);
assign soc_videooverlaysoc_core_mac_ps_crc_error_o = (soc_videooverlaysoc_core_mac_ps_crc_error_toggle_o ^ soc_videooverlaysoc_core_mac_ps_crc_error_toggle_o_r);
assign soc_videooverlaysoc_core_mac_padding_inserter_counter_done = (soc_videooverlaysoc_core_mac_padding_inserter_counter >= 6'd59);
always @(*) begin
	vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_next_state <= 1'd0;
	soc_videooverlaysoc_core_mac_padding_inserter_source_first <= 1'd0;
	soc_videooverlaysoc_core_mac_padding_inserter_source_last <= 1'd0;
	soc_videooverlaysoc_core_mac_padding_inserter_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_mac_padding_inserter_source_payload_last_be <= 1'd0;
	soc_videooverlaysoc_core_mac_padding_inserter_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_mac_padding_inserter_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_mac_padding_inserter_counter_ce <= 1'd0;
	soc_videooverlaysoc_core_mac_padding_inserter_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_mac_padding_inserter_source_valid <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_next_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_state;
	case (vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_state)
		1'd1: begin
			soc_videooverlaysoc_core_mac_padding_inserter_source_valid <= 1'd1;
			soc_videooverlaysoc_core_mac_padding_inserter_source_last <= soc_videooverlaysoc_core_mac_padding_inserter_counter_done;
			soc_videooverlaysoc_core_mac_padding_inserter_source_payload_data <= 1'd0;
			if ((soc_videooverlaysoc_core_mac_padding_inserter_source_valid & soc_videooverlaysoc_core_mac_padding_inserter_source_ready)) begin
				soc_videooverlaysoc_core_mac_padding_inserter_counter_ce <= 1'd1;
				if (soc_videooverlaysoc_core_mac_padding_inserter_counter_done) begin
					soc_videooverlaysoc_core_mac_padding_inserter_counter_reset <= 1'd1;
					vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_core_mac_padding_inserter_source_valid <= soc_videooverlaysoc_core_mac_padding_inserter_sink_valid;
			soc_videooverlaysoc_core_mac_padding_inserter_sink_ready <= soc_videooverlaysoc_core_mac_padding_inserter_source_ready;
			soc_videooverlaysoc_core_mac_padding_inserter_source_first <= soc_videooverlaysoc_core_mac_padding_inserter_sink_first;
			soc_videooverlaysoc_core_mac_padding_inserter_source_last <= soc_videooverlaysoc_core_mac_padding_inserter_sink_last;
			soc_videooverlaysoc_core_mac_padding_inserter_source_payload_data <= soc_videooverlaysoc_core_mac_padding_inserter_sink_payload_data;
			soc_videooverlaysoc_core_mac_padding_inserter_source_payload_last_be <= soc_videooverlaysoc_core_mac_padding_inserter_sink_payload_last_be;
			soc_videooverlaysoc_core_mac_padding_inserter_source_payload_error <= soc_videooverlaysoc_core_mac_padding_inserter_sink_payload_error;
			if ((soc_videooverlaysoc_core_mac_padding_inserter_source_valid & soc_videooverlaysoc_core_mac_padding_inserter_source_ready)) begin
				soc_videooverlaysoc_core_mac_padding_inserter_counter_ce <= 1'd1;
				if (soc_videooverlaysoc_core_mac_padding_inserter_sink_last) begin
					if ((~soc_videooverlaysoc_core_mac_padding_inserter_counter_done)) begin
						soc_videooverlaysoc_core_mac_padding_inserter_source_last <= 1'd0;
						vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_next_state <= 1'd1;
					end else begin
						soc_videooverlaysoc_core_mac_padding_inserter_counter_reset <= 1'd1;
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_mac_padding_checker_source_valid = soc_videooverlaysoc_core_mac_padding_checker_sink_valid;
assign soc_videooverlaysoc_core_mac_padding_checker_sink_ready = soc_videooverlaysoc_core_mac_padding_checker_source_ready;
assign soc_videooverlaysoc_core_mac_padding_checker_source_first = soc_videooverlaysoc_core_mac_padding_checker_sink_first;
assign soc_videooverlaysoc_core_mac_padding_checker_source_last = soc_videooverlaysoc_core_mac_padding_checker_sink_last;
assign soc_videooverlaysoc_core_mac_padding_checker_source_payload_data = soc_videooverlaysoc_core_mac_padding_checker_sink_payload_data;
assign soc_videooverlaysoc_core_mac_padding_checker_source_payload_last_be = soc_videooverlaysoc_core_mac_padding_checker_sink_payload_last_be;
assign soc_videooverlaysoc_core_mac_padding_checker_source_payload_error = soc_videooverlaysoc_core_mac_padding_checker_sink_payload_error;
assign soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_din = {soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_last, soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_first, soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_payload_error, soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_payload_last_be, soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_payload_data};
assign {soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_last, soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_first, soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_payload_error, soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_payload_last_be, soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_payload_data} = soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_dout;
assign soc_videooverlaysoc_core_mac_tx_cdc_sink_ready = soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_writable;
assign soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_we = soc_videooverlaysoc_core_mac_tx_cdc_sink_valid;
assign soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_first = soc_videooverlaysoc_core_mac_tx_cdc_sink_first;
assign soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_last = soc_videooverlaysoc_core_mac_tx_cdc_sink_last;
assign soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_payload_data = soc_videooverlaysoc_core_mac_tx_cdc_sink_payload_data;
assign soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_payload_last_be = soc_videooverlaysoc_core_mac_tx_cdc_sink_payload_last_be;
assign soc_videooverlaysoc_core_mac_tx_cdc_fifo_in_payload_error = soc_videooverlaysoc_core_mac_tx_cdc_sink_payload_error;
assign soc_videooverlaysoc_core_mac_tx_cdc_source_valid = soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_readable;
assign soc_videooverlaysoc_core_mac_tx_cdc_source_first = soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_first;
assign soc_videooverlaysoc_core_mac_tx_cdc_source_last = soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_last;
assign soc_videooverlaysoc_core_mac_tx_cdc_source_payload_data = soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_payload_data;
assign soc_videooverlaysoc_core_mac_tx_cdc_source_payload_last_be = soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_payload_last_be;
assign soc_videooverlaysoc_core_mac_tx_cdc_source_payload_error = soc_videooverlaysoc_core_mac_tx_cdc_fifo_out_payload_error;
assign soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_re = soc_videooverlaysoc_core_mac_tx_cdc_source_ready;
assign soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_ce = (soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_writable & soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_we);
assign soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_ce = (soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_readable & soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_re);
assign soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_writable = (((soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q[6] == soc_videooverlaysoc_core_mac_tx_cdc_consume_wdomain[6]) | (soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q[5] == soc_videooverlaysoc_core_mac_tx_cdc_consume_wdomain[5])) | (soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q[4:0] != soc_videooverlaysoc_core_mac_tx_cdc_consume_wdomain[4:0]));
assign soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_readable = (soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q != soc_videooverlaysoc_core_mac_tx_cdc_produce_rdomain);
assign soc_videooverlaysoc_core_mac_tx_cdc_wrport_adr = soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_binary[5:0];
assign soc_videooverlaysoc_core_mac_tx_cdc_wrport_dat_w = soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_din;
assign soc_videooverlaysoc_core_mac_tx_cdc_wrport_we = soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_ce;
assign soc_videooverlaysoc_core_mac_tx_cdc_rdport_adr = soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next_binary[5:0];
assign soc_videooverlaysoc_core_mac_tx_cdc_asyncfifo_dout = soc_videooverlaysoc_core_mac_tx_cdc_rdport_dat_r;
always @(*) begin
	soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_ce) begin
		soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_next_binary <= (soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_next_binary <= soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_binary;
	end
end
assign soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_next = (soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_next_binary ^ soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_next_binary[6:1]);
always @(*) begin
	soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_ce) begin
		soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next_binary <= (soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next_binary <= soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_binary;
	end
end
assign soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next = (soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next_binary ^ soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next_binary[6:1]);
assign soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_din = {soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_last, soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_first, soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_payload_error, soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_payload_last_be, soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_payload_data};
assign {soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_last, soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_first, soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_payload_error, soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_payload_last_be, soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_payload_data} = soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_dout;
assign soc_videooverlaysoc_core_mac_rx_cdc_sink_ready = soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_writable;
assign soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_we = soc_videooverlaysoc_core_mac_rx_cdc_sink_valid;
assign soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_first = soc_videooverlaysoc_core_mac_rx_cdc_sink_first;
assign soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_last = soc_videooverlaysoc_core_mac_rx_cdc_sink_last;
assign soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_payload_data = soc_videooverlaysoc_core_mac_rx_cdc_sink_payload_data;
assign soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_payload_last_be = soc_videooverlaysoc_core_mac_rx_cdc_sink_payload_last_be;
assign soc_videooverlaysoc_core_mac_rx_cdc_fifo_in_payload_error = soc_videooverlaysoc_core_mac_rx_cdc_sink_payload_error;
assign soc_videooverlaysoc_core_mac_rx_cdc_source_valid = soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_readable;
assign soc_videooverlaysoc_core_mac_rx_cdc_source_first = soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_first;
assign soc_videooverlaysoc_core_mac_rx_cdc_source_last = soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_last;
assign soc_videooverlaysoc_core_mac_rx_cdc_source_payload_data = soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_payload_data;
assign soc_videooverlaysoc_core_mac_rx_cdc_source_payload_last_be = soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_payload_last_be;
assign soc_videooverlaysoc_core_mac_rx_cdc_source_payload_error = soc_videooverlaysoc_core_mac_rx_cdc_fifo_out_payload_error;
assign soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_re = soc_videooverlaysoc_core_mac_rx_cdc_source_ready;
assign soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_ce = (soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_writable & soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_we);
assign soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_ce = (soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_readable & soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_re);
assign soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_writable = (((soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q[6] == soc_videooverlaysoc_core_mac_rx_cdc_consume_wdomain[6]) | (soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q[5] == soc_videooverlaysoc_core_mac_rx_cdc_consume_wdomain[5])) | (soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q[4:0] != soc_videooverlaysoc_core_mac_rx_cdc_consume_wdomain[4:0]));
assign soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_readable = (soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q != soc_videooverlaysoc_core_mac_rx_cdc_produce_rdomain);
assign soc_videooverlaysoc_core_mac_rx_cdc_wrport_adr = soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_binary[5:0];
assign soc_videooverlaysoc_core_mac_rx_cdc_wrport_dat_w = soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_din;
assign soc_videooverlaysoc_core_mac_rx_cdc_wrport_we = soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_ce;
assign soc_videooverlaysoc_core_mac_rx_cdc_rdport_adr = soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next_binary[5:0];
assign soc_videooverlaysoc_core_mac_rx_cdc_asyncfifo_dout = soc_videooverlaysoc_core_mac_rx_cdc_rdport_dat_r;
always @(*) begin
	soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_ce) begin
		soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_next_binary <= (soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_next_binary <= soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_binary;
	end
end
assign soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_next = (soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_next_binary ^ soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_next_binary[6:1]);
always @(*) begin
	soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_ce) begin
		soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next_binary <= (soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next_binary <= soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_binary;
	end
end
assign soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next = (soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next_binary ^ soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next_binary[6:1]);
assign soc_videooverlaysoc_core_mac_padding_inserter_sink_valid = soc_videooverlaysoc_core_mac_tx_cdc_source_valid;
assign soc_videooverlaysoc_core_mac_tx_cdc_source_ready = soc_videooverlaysoc_core_mac_padding_inserter_sink_ready;
assign soc_videooverlaysoc_core_mac_padding_inserter_sink_first = soc_videooverlaysoc_core_mac_tx_cdc_source_first;
assign soc_videooverlaysoc_core_mac_padding_inserter_sink_last = soc_videooverlaysoc_core_mac_tx_cdc_source_last;
assign soc_videooverlaysoc_core_mac_padding_inserter_sink_payload_data = soc_videooverlaysoc_core_mac_tx_cdc_source_payload_data;
assign soc_videooverlaysoc_core_mac_padding_inserter_sink_payload_last_be = soc_videooverlaysoc_core_mac_tx_cdc_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_padding_inserter_sink_payload_error = soc_videooverlaysoc_core_mac_tx_cdc_source_payload_error;
assign soc_videooverlaysoc_core_mac_crc32_inserter_sink_valid = soc_videooverlaysoc_core_mac_padding_inserter_source_valid;
assign soc_videooverlaysoc_core_mac_padding_inserter_source_ready = soc_videooverlaysoc_core_mac_crc32_inserter_sink_ready;
assign soc_videooverlaysoc_core_mac_crc32_inserter_sink_first = soc_videooverlaysoc_core_mac_padding_inserter_source_first;
assign soc_videooverlaysoc_core_mac_crc32_inserter_sink_last = soc_videooverlaysoc_core_mac_padding_inserter_source_last;
assign soc_videooverlaysoc_core_mac_crc32_inserter_sink_payload_data = soc_videooverlaysoc_core_mac_padding_inserter_source_payload_data;
assign soc_videooverlaysoc_core_mac_crc32_inserter_sink_payload_last_be = soc_videooverlaysoc_core_mac_padding_inserter_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_crc32_inserter_sink_payload_error = soc_videooverlaysoc_core_mac_padding_inserter_source_payload_error;
assign soc_videooverlaysoc_core_mac_preamble_inserter_sink_valid = soc_videooverlaysoc_core_mac_crc32_inserter_source_valid;
assign soc_videooverlaysoc_core_mac_crc32_inserter_source_ready = soc_videooverlaysoc_core_mac_preamble_inserter_sink_ready;
assign soc_videooverlaysoc_core_mac_preamble_inserter_sink_first = soc_videooverlaysoc_core_mac_crc32_inserter_source_first;
assign soc_videooverlaysoc_core_mac_preamble_inserter_sink_last = soc_videooverlaysoc_core_mac_crc32_inserter_source_last;
assign soc_videooverlaysoc_core_mac_preamble_inserter_sink_payload_data = soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_data;
assign soc_videooverlaysoc_core_mac_preamble_inserter_sink_payload_last_be = soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_preamble_inserter_sink_payload_error = soc_videooverlaysoc_core_mac_crc32_inserter_source_payload_error;
assign soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_valid = soc_videooverlaysoc_core_mac_preamble_inserter_source_valid;
assign soc_videooverlaysoc_core_mac_preamble_inserter_source_ready = soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_ready;
assign soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_first = soc_videooverlaysoc_core_mac_preamble_inserter_source_first;
assign soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_last = soc_videooverlaysoc_core_mac_preamble_inserter_source_last;
assign soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_payload_data = soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_data;
assign soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_payload_last_be = soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_tx_gap_inserter_sink_payload_error = soc_videooverlaysoc_core_mac_preamble_inserter_source_payload_error;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_valid = soc_videooverlaysoc_core_mac_tx_gap_inserter_source_valid;
assign soc_videooverlaysoc_core_mac_tx_gap_inserter_source_ready = soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_ready;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_first = soc_videooverlaysoc_core_mac_tx_gap_inserter_source_first;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_last = soc_videooverlaysoc_core_mac_tx_gap_inserter_source_last;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_payload_data = soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_data;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_payload_last_be = soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_last_be;
assign soc_videooverlaysoc_phy_liteethphyrmiitx_sink_sink_payload_error = soc_videooverlaysoc_core_mac_tx_gap_inserter_source_payload_error;
assign soc_videooverlaysoc_core_mac_preamble_checker_sink_valid = soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_valid;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_ready = soc_videooverlaysoc_core_mac_preamble_checker_sink_ready;
assign soc_videooverlaysoc_core_mac_preamble_checker_sink_first = soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_first;
assign soc_videooverlaysoc_core_mac_preamble_checker_sink_last = soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_last;
assign soc_videooverlaysoc_core_mac_preamble_checker_sink_payload_data = soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_payload_data;
assign soc_videooverlaysoc_core_mac_preamble_checker_sink_payload_last_be = soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_preamble_checker_sink_payload_error = soc_videooverlaysoc_phy_liteethphyrmiirx_source_source_payload_error;
assign soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_valid = soc_videooverlaysoc_core_mac_preamble_checker_source_valid;
assign soc_videooverlaysoc_core_mac_preamble_checker_source_ready = soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_ready;
assign soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_first = soc_videooverlaysoc_core_mac_preamble_checker_source_first;
assign soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_last = soc_videooverlaysoc_core_mac_preamble_checker_source_last;
assign soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_data = soc_videooverlaysoc_core_mac_preamble_checker_source_payload_data;
assign soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_last_be = soc_videooverlaysoc_core_mac_preamble_checker_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_crc32_checker_sink_sink_payload_error = soc_videooverlaysoc_core_mac_preamble_checker_source_payload_error;
assign soc_videooverlaysoc_core_mac_padding_checker_sink_valid = soc_videooverlaysoc_core_mac_crc32_checker_source_source_valid;
assign soc_videooverlaysoc_core_mac_crc32_checker_source_source_ready = soc_videooverlaysoc_core_mac_padding_checker_sink_ready;
assign soc_videooverlaysoc_core_mac_padding_checker_sink_first = soc_videooverlaysoc_core_mac_crc32_checker_source_source_first;
assign soc_videooverlaysoc_core_mac_padding_checker_sink_last = soc_videooverlaysoc_core_mac_crc32_checker_source_source_last;
assign soc_videooverlaysoc_core_mac_padding_checker_sink_payload_data = soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_data;
assign soc_videooverlaysoc_core_mac_padding_checker_sink_payload_last_be = soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_padding_checker_sink_payload_error = soc_videooverlaysoc_core_mac_crc32_checker_source_source_payload_error;
assign soc_videooverlaysoc_core_mac_rx_cdc_sink_valid = soc_videooverlaysoc_core_mac_padding_checker_source_valid;
assign soc_videooverlaysoc_core_mac_padding_checker_source_ready = soc_videooverlaysoc_core_mac_rx_cdc_sink_ready;
assign soc_videooverlaysoc_core_mac_rx_cdc_sink_first = soc_videooverlaysoc_core_mac_padding_checker_source_first;
assign soc_videooverlaysoc_core_mac_rx_cdc_sink_last = soc_videooverlaysoc_core_mac_padding_checker_source_last;
assign soc_videooverlaysoc_core_mac_rx_cdc_sink_payload_data = soc_videooverlaysoc_core_mac_padding_checker_source_payload_data;
assign soc_videooverlaysoc_core_mac_rx_cdc_sink_payload_last_be = soc_videooverlaysoc_core_mac_padding_checker_source_payload_last_be;
assign soc_videooverlaysoc_core_mac_rx_cdc_sink_payload_error = soc_videooverlaysoc_core_mac_padding_checker_source_payload_error;
always @(*) begin
	vns_clockdomainsrenamer1_liteethmac_sel0 <= 2'd0;
	case (soc_videooverlaysoc_core_mac_crossbar_sink_payload_ethernet_type)
		12'd2048: begin
			vns_clockdomainsrenamer1_liteethmac_sel0 <= 2'd2;
		end
		12'd2054: begin
			vns_clockdomainsrenamer1_liteethmac_sel0 <= 1'd1;
		end
		default: begin
			vns_clockdomainsrenamer1_liteethmac_sel0 <= 1'd0;
		end
	endcase
end
always @(*) begin
	vns_clockdomainsrenamer1_liteethmac_request <= 2'd0;
	vns_clockdomainsrenamer1_liteethmac_request[0] <= vns_clockdomainsrenamer1_liteethmac_status0_ongoing0;
	vns_clockdomainsrenamer1_liteethmac_request[1] <= vns_clockdomainsrenamer1_liteethmac_status1_ongoing0;
end
always @(*) begin
	soc_videooverlaysoc_core_mac_crossbar_source_valid <= 1'd0;
	soc_videooverlaysoc_core_mac_crossbar_source_first <= 1'd0;
	soc_videooverlaysoc_core_mac_crossbar_source_last <= 1'd0;
	soc_videooverlaysoc_core_mac_crossbar_source_payload_ethernet_type <= 16'd0;
	soc_videooverlaysoc_core_mac_crossbar_source_payload_sender_mac <= 48'd0;
	soc_videooverlaysoc_core_mac_crossbar_source_payload_target_mac <= 48'd0;
	soc_videooverlaysoc_core_mac_crossbar_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_mac_crossbar_source_payload_last_be <= 1'd0;
	soc_videooverlaysoc_core_mac_crossbar_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_arp_mac_port_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_ip_mac_port_sink_ready <= 1'd0;
	case (vns_clockdomainsrenamer1_liteethmac_grant)
		1'd0: begin
			soc_videooverlaysoc_core_mac_crossbar_source_valid <= soc_videooverlaysoc_core_arp_mac_port_sink_valid;
			soc_videooverlaysoc_core_arp_mac_port_sink_ready <= soc_videooverlaysoc_core_mac_crossbar_source_ready;
			soc_videooverlaysoc_core_mac_crossbar_source_first <= soc_videooverlaysoc_core_arp_mac_port_sink_first;
			soc_videooverlaysoc_core_mac_crossbar_source_last <= soc_videooverlaysoc_core_arp_mac_port_sink_last;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_ethernet_type <= soc_videooverlaysoc_core_arp_mac_port_sink_payload_ethernet_type;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_sender_mac <= soc_videooverlaysoc_core_arp_mac_port_sink_payload_sender_mac;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_target_mac <= soc_videooverlaysoc_core_arp_mac_port_sink_payload_target_mac;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_data <= soc_videooverlaysoc_core_arp_mac_port_sink_payload_data;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_last_be <= soc_videooverlaysoc_core_arp_mac_port_sink_payload_last_be;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_error <= soc_videooverlaysoc_core_arp_mac_port_sink_payload_error;
		end
		1'd1: begin
			soc_videooverlaysoc_core_mac_crossbar_source_valid <= soc_videooverlaysoc_core_ip_mac_port_sink_valid;
			soc_videooverlaysoc_core_ip_mac_port_sink_ready <= soc_videooverlaysoc_core_mac_crossbar_source_ready;
			soc_videooverlaysoc_core_mac_crossbar_source_first <= soc_videooverlaysoc_core_ip_mac_port_sink_first;
			soc_videooverlaysoc_core_mac_crossbar_source_last <= soc_videooverlaysoc_core_ip_mac_port_sink_last;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_ethernet_type <= soc_videooverlaysoc_core_ip_mac_port_sink_payload_ethernet_type;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_sender_mac <= soc_videooverlaysoc_core_ip_mac_port_sink_payload_sender_mac;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_target_mac <= soc_videooverlaysoc_core_ip_mac_port_sink_payload_target_mac;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_data <= soc_videooverlaysoc_core_ip_mac_port_sink_payload_data;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_last_be <= soc_videooverlaysoc_core_ip_mac_port_sink_payload_last_be;
			soc_videooverlaysoc_core_mac_crossbar_source_payload_error <= soc_videooverlaysoc_core_ip_mac_port_sink_payload_error;
		end
	endcase
end
always @(*) begin
	vns_clockdomainsrenamer1_liteethmac_status0_last <= 1'd0;
	if (soc_videooverlaysoc_core_arp_mac_port_sink_valid) begin
		vns_clockdomainsrenamer1_liteethmac_status0_last <= (soc_videooverlaysoc_core_arp_mac_port_sink_last & soc_videooverlaysoc_core_arp_mac_port_sink_ready);
	end
end
assign vns_clockdomainsrenamer1_liteethmac_status0_ongoing0 = ((soc_videooverlaysoc_core_arp_mac_port_sink_valid | vns_clockdomainsrenamer1_liteethmac_status0_ongoing1) & (~vns_clockdomainsrenamer1_liteethmac_status0_last));
always @(*) begin
	vns_clockdomainsrenamer1_liteethmac_status1_last <= 1'd0;
	if (soc_videooverlaysoc_core_ip_mac_port_sink_valid) begin
		vns_clockdomainsrenamer1_liteethmac_status1_last <= (soc_videooverlaysoc_core_ip_mac_port_sink_last & soc_videooverlaysoc_core_ip_mac_port_sink_ready);
	end
end
assign vns_clockdomainsrenamer1_liteethmac_status1_ongoing0 = ((soc_videooverlaysoc_core_ip_mac_port_sink_valid | vns_clockdomainsrenamer1_liteethmac_status1_ongoing1) & (~vns_clockdomainsrenamer1_liteethmac_status1_last));
always @(*) begin
	vns_clockdomainsrenamer1_liteethmac_sel1 <= 2'd0;
	if (vns_clockdomainsrenamer1_liteethmac_first) begin
		vns_clockdomainsrenamer1_liteethmac_sel1 <= vns_clockdomainsrenamer1_liteethmac_sel0;
	end else begin
		vns_clockdomainsrenamer1_liteethmac_sel1 <= vns_clockdomainsrenamer1_liteethmac_sel_ongoing;
	end
end
always @(*) begin
	soc_videooverlaysoc_core_arp_mac_port_source_valid <= 1'd0;
	soc_videooverlaysoc_core_arp_mac_port_source_first <= 1'd0;
	soc_videooverlaysoc_core_arp_mac_port_source_last <= 1'd0;
	soc_videooverlaysoc_core_arp_mac_port_source_payload_ethernet_type <= 16'd0;
	soc_videooverlaysoc_core_arp_mac_port_source_payload_sender_mac <= 48'd0;
	soc_videooverlaysoc_core_ip_mac_port_source_valid <= 1'd0;
	soc_videooverlaysoc_core_arp_mac_port_source_payload_target_mac <= 48'd0;
	soc_videooverlaysoc_core_arp_mac_port_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_ip_mac_port_source_first <= 1'd0;
	soc_videooverlaysoc_core_arp_mac_port_source_payload_last_be <= 1'd0;
	soc_videooverlaysoc_core_mac_crossbar_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_ip_mac_port_source_payload_ethernet_type <= 16'd0;
	soc_videooverlaysoc_core_arp_mac_port_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_ip_mac_port_source_last <= 1'd0;
	soc_videooverlaysoc_core_ip_mac_port_source_payload_sender_mac <= 48'd0;
	soc_videooverlaysoc_core_ip_mac_port_source_payload_target_mac <= 48'd0;
	soc_videooverlaysoc_core_ip_mac_port_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_ip_mac_port_source_payload_last_be <= 1'd0;
	soc_videooverlaysoc_core_ip_mac_port_source_payload_error <= 1'd0;
	case (vns_clockdomainsrenamer1_liteethmac_sel1)
		1'd1: begin
			soc_videooverlaysoc_core_arp_mac_port_source_valid <= soc_videooverlaysoc_core_mac_crossbar_sink_valid;
			soc_videooverlaysoc_core_mac_crossbar_sink_ready <= soc_videooverlaysoc_core_arp_mac_port_source_ready;
			soc_videooverlaysoc_core_arp_mac_port_source_first <= soc_videooverlaysoc_core_mac_crossbar_sink_first;
			soc_videooverlaysoc_core_arp_mac_port_source_last <= soc_videooverlaysoc_core_mac_crossbar_sink_last;
			soc_videooverlaysoc_core_arp_mac_port_source_payload_ethernet_type <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_ethernet_type;
			soc_videooverlaysoc_core_arp_mac_port_source_payload_sender_mac <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_sender_mac;
			soc_videooverlaysoc_core_arp_mac_port_source_payload_target_mac <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_target_mac;
			soc_videooverlaysoc_core_arp_mac_port_source_payload_data <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_data;
			soc_videooverlaysoc_core_arp_mac_port_source_payload_last_be <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_last_be;
			soc_videooverlaysoc_core_arp_mac_port_source_payload_error <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_error;
		end
		2'd2: begin
			soc_videooverlaysoc_core_ip_mac_port_source_valid <= soc_videooverlaysoc_core_mac_crossbar_sink_valid;
			soc_videooverlaysoc_core_mac_crossbar_sink_ready <= soc_videooverlaysoc_core_ip_mac_port_source_ready;
			soc_videooverlaysoc_core_ip_mac_port_source_first <= soc_videooverlaysoc_core_mac_crossbar_sink_first;
			soc_videooverlaysoc_core_ip_mac_port_source_last <= soc_videooverlaysoc_core_mac_crossbar_sink_last;
			soc_videooverlaysoc_core_ip_mac_port_source_payload_ethernet_type <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_ethernet_type;
			soc_videooverlaysoc_core_ip_mac_port_source_payload_sender_mac <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_sender_mac;
			soc_videooverlaysoc_core_ip_mac_port_source_payload_target_mac <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_target_mac;
			soc_videooverlaysoc_core_ip_mac_port_source_payload_data <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_data;
			soc_videooverlaysoc_core_ip_mac_port_source_payload_last_be <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_last_be;
			soc_videooverlaysoc_core_ip_mac_port_source_payload_error <= soc_videooverlaysoc_core_mac_crossbar_sink_payload_error;
		end
		default: begin
			soc_videooverlaysoc_core_mac_crossbar_sink_ready <= 1'd1;
		end
	endcase
end
always @(*) begin
	vns_clockdomainsrenamer1_liteethmac_last <= 1'd0;
	if (soc_videooverlaysoc_core_mac_crossbar_sink_valid) begin
		vns_clockdomainsrenamer1_liteethmac_last <= (soc_videooverlaysoc_core_mac_crossbar_sink_last & soc_videooverlaysoc_core_mac_crossbar_sink_ready);
	end
end
assign vns_clockdomainsrenamer1_liteethmac_ongoing0 = ((soc_videooverlaysoc_core_mac_crossbar_sink_valid | vns_clockdomainsrenamer1_liteethmac_ongoing1) & (~vns_clockdomainsrenamer1_liteethmac_last));
always @(*) begin
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_header <= 112'd0;
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_header[111:96] <= {soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_ethernet_type[7:0], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_ethernet_type[15:8]};
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_header[95:48] <= {soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_sender_mac[7:0], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_sender_mac[15:8], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_sender_mac[23:16], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_sender_mac[31:24], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_sender_mac[39:32], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_sender_mac[47:40]};
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_header[47:0] <= {soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_target_mac[7:0], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_target_mac[15:8], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_target_mac[23:16], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_target_mac[31:24], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_target_mac[39:32], soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_target_mac[47:40]};
end
assign soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_error = soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_error;
always @(*) begin
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_last <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_next_state <= 2'd0;
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_load <= 1'd0;
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_shift <= 1'd0;
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter_ce <= 1'd0;
	soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_valid <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_next_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_state;
	case (vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_valid <= 1'd1;
			soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_last <= 1'd0;
			soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_data <= soc_videooverlaysoc_core_mac_liteethmacpacketizer_header_reg[15:8];
			if ((soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_valid & soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_ready)) begin
				soc_videooverlaysoc_core_mac_liteethmacpacketizer_shift <= 1'd1;
				soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter_ce <= 1'd1;
				if ((soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter == 4'd12)) begin
					vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_valid <= soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_valid;
			soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_last <= soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_last;
			soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_data <= soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_payload_data;
			if ((soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_valid & soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_ready)) begin
				soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_ready <= 1'd1;
				if (soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_last) begin
					vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_valid) begin
				soc_videooverlaysoc_core_mac_liteethmacpacketizer_sink_ready <= 1'd0;
				soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_valid <= 1'd1;
				soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_last <= 1'd0;
				soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_payload_data <= soc_videooverlaysoc_core_mac_liteethmacpacketizer_header[7:0];
				if ((soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_valid & soc_videooverlaysoc_core_mac_liteethmacpacketizer_source_ready)) begin
					soc_videooverlaysoc_core_mac_liteethmacpacketizer_load <= 1'd1;
					vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_next_state <= 1'd1;
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_mac_depacketizer_header = soc_videooverlaysoc_core_mac_depacketizer_header_reg;
assign soc_videooverlaysoc_core_mac_depacketizer_source_payload_error = soc_videooverlaysoc_core_mac_depacketizer_sink_payload_error;
assign soc_videooverlaysoc_core_mac_depacketizer_source_last = (soc_videooverlaysoc_core_mac_depacketizer_sink_last | soc_videooverlaysoc_core_mac_depacketizer_no_payload);
assign soc_videooverlaysoc_core_mac_depacketizer_source_payload_data = soc_videooverlaysoc_core_mac_depacketizer_sink_payload_data;
assign soc_videooverlaysoc_core_mac_depacketizer_source_payload_ethernet_type = {vns_slice_proxy1[7:0], vns_slice_proxy0[15:8]};
assign soc_videooverlaysoc_core_mac_depacketizer_source_payload_sender_mac = {vns_slice_proxy7[7:0], vns_slice_proxy6[15:8], vns_slice_proxy5[23:16], vns_slice_proxy4[31:24], vns_slice_proxy3[39:32], vns_slice_proxy2[47:40]};
assign soc_videooverlaysoc_core_mac_depacketizer_source_payload_target_mac = {vns_slice_proxy13[7:0], vns_slice_proxy12[15:8], vns_slice_proxy11[23:16], vns_slice_proxy10[31:24], vns_slice_proxy9[39:32], vns_slice_proxy8[47:40]};
always @(*) begin
	soc_videooverlaysoc_core_mac_depacketizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_mac_depacketizer_counter_ce <= 1'd0;
	soc_videooverlaysoc_core_mac_depacketizer_source_valid <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_next_state <= 2'd0;
	soc_videooverlaysoc_core_mac_depacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_mac_depacketizer_shift <= 1'd0;
	vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_next_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_state;
	case (vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_core_mac_depacketizer_sink_ready <= 1'd1;
			if (soc_videooverlaysoc_core_mac_depacketizer_sink_valid) begin
				soc_videooverlaysoc_core_mac_depacketizer_counter_ce <= 1'd1;
				soc_videooverlaysoc_core_mac_depacketizer_shift <= 1'd1;
				if ((soc_videooverlaysoc_core_mac_depacketizer_counter == 4'd12)) begin
					vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_mac_depacketizer_sink_ready <= soc_videooverlaysoc_core_mac_depacketizer_source_ready;
			soc_videooverlaysoc_core_mac_depacketizer_source_valid <= (soc_videooverlaysoc_core_mac_depacketizer_sink_valid | soc_videooverlaysoc_core_mac_depacketizer_no_payload);
			if (((soc_videooverlaysoc_core_mac_depacketizer_source_valid & soc_videooverlaysoc_core_mac_depacketizer_source_ready) & soc_videooverlaysoc_core_mac_depacketizer_source_last)) begin
				vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_mac_depacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_mac_depacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_mac_depacketizer_sink_valid) begin
				soc_videooverlaysoc_core_mac_depacketizer_shift <= 1'd1;
				vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_mac_depacketizer_is_el = ((~(vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_state == 2'd2)) & (vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_next_state == 2'd2));
assign soc_videooverlaysoc_core_arp_table_sink_valid = soc_videooverlaysoc_core_arp_source_source_valid;
assign soc_videooverlaysoc_core_arp_source_source_ready = soc_videooverlaysoc_core_arp_table_sink_ready;
assign soc_videooverlaysoc_core_arp_table_sink_first = soc_videooverlaysoc_core_arp_source_source_first;
assign soc_videooverlaysoc_core_arp_table_sink_last = soc_videooverlaysoc_core_arp_source_source_last;
assign soc_videooverlaysoc_core_arp_table_sink_payload_reply = soc_videooverlaysoc_core_arp_source_source_payload_reply;
assign soc_videooverlaysoc_core_arp_table_sink_payload_request = soc_videooverlaysoc_core_arp_source_source_payload_request;
assign soc_videooverlaysoc_core_arp_table_sink_payload_ip_address = soc_videooverlaysoc_core_arp_source_source_payload_ip_address;
assign soc_videooverlaysoc_core_arp_table_sink_payload_mac_address = soc_videooverlaysoc_core_arp_source_source_payload_mac_address;
assign soc_videooverlaysoc_core_arp_tx_sink_valid = soc_videooverlaysoc_core_arp_table_source_valid;
assign soc_videooverlaysoc_core_arp_table_source_ready = soc_videooverlaysoc_core_arp_tx_sink_ready;
assign soc_videooverlaysoc_core_arp_tx_sink_first = soc_videooverlaysoc_core_arp_table_source_first;
assign soc_videooverlaysoc_core_arp_tx_sink_last = soc_videooverlaysoc_core_arp_table_source_last;
assign soc_videooverlaysoc_core_arp_tx_sink_payload_reply = soc_videooverlaysoc_core_arp_table_source_payload_reply;
assign soc_videooverlaysoc_core_arp_tx_sink_payload_request = soc_videooverlaysoc_core_arp_table_source_payload_request;
assign soc_videooverlaysoc_core_arp_tx_sink_payload_ip_address = soc_videooverlaysoc_core_arp_table_source_payload_ip_address;
assign soc_videooverlaysoc_core_arp_tx_sink_payload_mac_address = soc_videooverlaysoc_core_arp_table_source_payload_mac_address;
assign soc_videooverlaysoc_core_arp_mac_port_sink_valid = soc_videooverlaysoc_core_arp_tx_source_valid;
assign soc_videooverlaysoc_core_arp_tx_source_ready = soc_videooverlaysoc_core_arp_mac_port_sink_ready;
assign soc_videooverlaysoc_core_arp_mac_port_sink_first = soc_videooverlaysoc_core_arp_tx_source_first;
assign soc_videooverlaysoc_core_arp_mac_port_sink_last = soc_videooverlaysoc_core_arp_tx_source_last;
assign soc_videooverlaysoc_core_arp_mac_port_sink_payload_ethernet_type = soc_videooverlaysoc_core_arp_tx_source_payload_ethernet_type;
assign soc_videooverlaysoc_core_arp_mac_port_sink_payload_sender_mac = soc_videooverlaysoc_core_arp_tx_source_payload_sender_mac;
assign soc_videooverlaysoc_core_arp_mac_port_sink_payload_target_mac = soc_videooverlaysoc_core_arp_tx_source_payload_target_mac;
assign soc_videooverlaysoc_core_arp_mac_port_sink_payload_data = soc_videooverlaysoc_core_arp_tx_source_payload_data;
assign soc_videooverlaysoc_core_arp_mac_port_sink_payload_last_be = soc_videooverlaysoc_core_arp_tx_source_payload_last_be;
assign soc_videooverlaysoc_core_arp_mac_port_sink_payload_error = soc_videooverlaysoc_core_arp_tx_source_payload_error;
assign soc_videooverlaysoc_core_arp_sink_sink_valid = soc_videooverlaysoc_core_arp_mac_port_source_valid;
assign soc_videooverlaysoc_core_arp_mac_port_source_ready = soc_videooverlaysoc_core_arp_sink_sink_ready;
assign soc_videooverlaysoc_core_arp_sink_sink_first = soc_videooverlaysoc_core_arp_mac_port_source_first;
assign soc_videooverlaysoc_core_arp_sink_sink_last = soc_videooverlaysoc_core_arp_mac_port_source_last;
assign soc_videooverlaysoc_core_arp_sink_sink_payload_ethernet_type = soc_videooverlaysoc_core_arp_mac_port_source_payload_ethernet_type;
assign soc_videooverlaysoc_core_arp_sink_sink_payload_sender_mac = soc_videooverlaysoc_core_arp_mac_port_source_payload_sender_mac;
assign soc_videooverlaysoc_core_arp_sink_sink_payload_target_mac = soc_videooverlaysoc_core_arp_mac_port_source_payload_target_mac;
assign soc_videooverlaysoc_core_arp_sink_sink_payload_data = soc_videooverlaysoc_core_arp_mac_port_source_payload_data;
assign soc_videooverlaysoc_core_arp_sink_sink_payload_last_be = soc_videooverlaysoc_core_arp_mac_port_source_payload_last_be;
assign soc_videooverlaysoc_core_arp_sink_sink_payload_error = soc_videooverlaysoc_core_arp_mac_port_source_payload_error;
assign soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_last = (soc_videooverlaysoc_core_arp_tx_counter == 6'd45);
assign soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_hwtype = 1'd1;
assign soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_proto = 12'd2048;
assign soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_hwsize = 3'd6;
assign soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_protosize = 3'd4;
assign soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_mac = 45'd21127783889598;
assign soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_ip = 28'd167774978;
always @(*) begin
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_opcode <= 16'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_ip <= 32'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac <= 48'd0;
	if (soc_videooverlaysoc_core_arp_tx_sink_payload_reply) begin
		soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_opcode <= 2'd2;
		soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac <= soc_videooverlaysoc_core_arp_tx_sink_payload_mac_address;
		soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_ip <= soc_videooverlaysoc_core_arp_tx_sink_payload_ip_address;
	end else begin
		if (soc_videooverlaysoc_core_arp_tx_sink_payload_request) begin
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_opcode <= 1'd1;
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac <= 48'd281474976710655;
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_ip <= soc_videooverlaysoc_core_arp_tx_sink_payload_ip_address;
		end
	end
end
always @(*) begin
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header <= 224'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header[39:32] <= {soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_hwsize[7:0]};
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header[15:0] <= {soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_hwtype[7:0], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_hwtype[15:8]};
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header[63:48] <= {soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_opcode[7:0], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_opcode[15:8]};
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header[31:16] <= {soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_proto[7:0], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_proto[15:8]};
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header[47:40] <= {soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_protosize[7:0]};
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header[143:112] <= {soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_ip[7:0], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_ip[15:8], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_ip[23:16], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_ip[31:24]};
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header[111:64] <= {soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_mac[7:0], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_mac[15:8], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_mac[23:16], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_mac[31:24], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_mac[39:32], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_sender_mac[47:40]};
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header[223:192] <= {soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_ip[7:0], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_ip[15:8], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_ip[23:16], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_ip[31:24]};
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header[191:144] <= {soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac[7:0], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac[15:8], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac[23:16], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac[31:24], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac[39:32], soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac[47:40]};
end
assign soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_error = soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_payload_error;
always @(*) begin
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_last <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_data <= 8'd0;
	vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_next_state <= 2'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_valid <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_load <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_shift <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter_ce <= 1'd0;
	vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_next_state <= vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_state;
	case (vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_valid <= 1'd1;
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_last <= 1'd0;
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_data <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header_reg[15:8];
			if ((soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_valid & soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_ready)) begin
				soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_shift <= 1'd1;
				soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter_ce <= 1'd1;
				if ((soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter == 5'd26)) begin
					vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_valid <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_valid;
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_last <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_last;
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_data <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_payload_data;
			if ((soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_valid & soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_ready)) begin
				soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_ready <= 1'd1;
				if (soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_last) begin
					vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_valid) begin
				soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_ready <= 1'd0;
				soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_valid <= 1'd1;
				soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_last <= 1'd0;
				soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_data <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header[7:0];
				if ((soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_valid & soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_ready)) begin
					soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_load <= 1'd1;
					vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_next_state <= 1'd1;
				end
			end
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_valid <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_ready <= 1'd0;
	vns_clockdomainsrenamer1_liteetharptx_fsm_next_state <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_counter_ce <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_source_valid <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_source_first <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_source_last <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_source_payload_ethernet_type <= 16'd0;
	soc_videooverlaysoc_core_arp_tx_source_payload_sender_mac <= 48'd0;
	soc_videooverlaysoc_core_arp_tx_source_payload_target_mac <= 48'd0;
	soc_videooverlaysoc_core_arp_tx_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_arp_tx_source_payload_last_be <= 1'd0;
	soc_videooverlaysoc_core_arp_tx_source_payload_error <= 1'd0;
	vns_clockdomainsrenamer1_liteetharptx_fsm_next_state <= vns_clockdomainsrenamer1_liteetharptx_fsm_state;
	case (vns_clockdomainsrenamer1_liteetharptx_fsm_state)
		1'd1: begin
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_valid <= 1'd1;
			soc_videooverlaysoc_core_arp_tx_source_valid <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_valid;
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_ready <= soc_videooverlaysoc_core_arp_tx_source_ready;
			soc_videooverlaysoc_core_arp_tx_source_first <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_first;
			soc_videooverlaysoc_core_arp_tx_source_last <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_last;
			soc_videooverlaysoc_core_arp_tx_source_payload_ethernet_type <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_ethernet_type;
			soc_videooverlaysoc_core_arp_tx_source_payload_sender_mac <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_sender_mac;
			soc_videooverlaysoc_core_arp_tx_source_payload_target_mac <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_target_mac;
			soc_videooverlaysoc_core_arp_tx_source_payload_data <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_data;
			soc_videooverlaysoc_core_arp_tx_source_payload_last_be <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_last_be;
			soc_videooverlaysoc_core_arp_tx_source_payload_error <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_source_payload_error;
			soc_videooverlaysoc_core_arp_tx_source_payload_target_mac <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_sink_param_target_mac;
			soc_videooverlaysoc_core_arp_tx_source_payload_sender_mac <= 45'd21127783889598;
			soc_videooverlaysoc_core_arp_tx_source_payload_ethernet_type <= 12'd2054;
			if ((soc_videooverlaysoc_core_arp_tx_source_valid & soc_videooverlaysoc_core_arp_tx_source_ready)) begin
				soc_videooverlaysoc_core_arp_tx_counter_ce <= 1'd1;
				if (soc_videooverlaysoc_core_arp_tx_source_last) begin
					soc_videooverlaysoc_core_arp_tx_sink_ready <= 1'd1;
					vns_clockdomainsrenamer1_liteetharptx_fsm_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_core_arp_tx_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_arp_tx_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_arp_tx_sink_valid) begin
				soc_videooverlaysoc_core_arp_tx_sink_ready <= 1'd0;
				vns_clockdomainsrenamer1_liteetharptx_fsm_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_arp_depacketizer_sink_valid = soc_videooverlaysoc_core_arp_sink_sink_valid;
assign soc_videooverlaysoc_core_arp_sink_sink_ready = soc_videooverlaysoc_core_arp_depacketizer_sink_ready;
assign soc_videooverlaysoc_core_arp_depacketizer_sink_first = soc_videooverlaysoc_core_arp_sink_sink_first;
assign soc_videooverlaysoc_core_arp_depacketizer_sink_last = soc_videooverlaysoc_core_arp_sink_sink_last;
assign soc_videooverlaysoc_core_arp_depacketizer_sink_payload_ethernet_type = soc_videooverlaysoc_core_arp_sink_sink_payload_ethernet_type;
assign soc_videooverlaysoc_core_arp_depacketizer_sink_payload_sender_mac = soc_videooverlaysoc_core_arp_sink_sink_payload_sender_mac;
assign soc_videooverlaysoc_core_arp_depacketizer_sink_payload_target_mac = soc_videooverlaysoc_core_arp_sink_sink_payload_target_mac;
assign soc_videooverlaysoc_core_arp_depacketizer_sink_payload_data = soc_videooverlaysoc_core_arp_sink_sink_payload_data;
assign soc_videooverlaysoc_core_arp_depacketizer_sink_payload_last_be = soc_videooverlaysoc_core_arp_sink_sink_payload_last_be;
assign soc_videooverlaysoc_core_arp_depacketizer_sink_payload_error = soc_videooverlaysoc_core_arp_sink_sink_payload_error;
always @(*) begin
	soc_videooverlaysoc_core_arp_reply <= 1'd0;
	soc_videooverlaysoc_core_arp_request <= 1'd0;
	case (soc_videooverlaysoc_core_arp_depacketizer_source_param_opcode)
		1'd1: begin
			soc_videooverlaysoc_core_arp_request <= 1'd1;
		end
		2'd2: begin
			soc_videooverlaysoc_core_arp_reply <= 1'd1;
		end
		default: begin
		end
	endcase
end
assign soc_videooverlaysoc_core_arp_source_source_payload_ip_address = soc_videooverlaysoc_core_arp_depacketizer_source_param_sender_ip;
assign soc_videooverlaysoc_core_arp_source_source_payload_mac_address = soc_videooverlaysoc_core_arp_depacketizer_source_param_sender_mac;
assign soc_videooverlaysoc_core_arp_depacketizer_header = soc_videooverlaysoc_core_arp_depacketizer_header_reg;
assign soc_videooverlaysoc_core_arp_depacketizer_source_payload_error = soc_videooverlaysoc_core_arp_depacketizer_sink_payload_error;
assign soc_videooverlaysoc_core_arp_depacketizer_source_last = (soc_videooverlaysoc_core_arp_depacketizer_sink_last | soc_videooverlaysoc_core_arp_depacketizer_no_payload);
assign soc_videooverlaysoc_core_arp_depacketizer_source_payload_data = soc_videooverlaysoc_core_arp_depacketizer_sink_payload_data;
assign soc_videooverlaysoc_core_arp_depacketizer_source_param_hwsize = {vns_slice_proxy14[7:0]};
assign soc_videooverlaysoc_core_arp_depacketizer_source_param_hwtype = {vns_slice_proxy16[7:0], vns_slice_proxy15[15:8]};
assign soc_videooverlaysoc_core_arp_depacketizer_source_param_opcode = {vns_slice_proxy18[7:0], vns_slice_proxy17[15:8]};
assign soc_videooverlaysoc_core_arp_depacketizer_source_param_proto = {vns_slice_proxy20[7:0], vns_slice_proxy19[15:8]};
assign soc_videooverlaysoc_core_arp_depacketizer_source_param_protosize = {vns_slice_proxy21[7:0]};
assign soc_videooverlaysoc_core_arp_depacketizer_source_param_sender_ip = {vns_slice_proxy25[7:0], vns_slice_proxy24[15:8], vns_slice_proxy23[23:16], vns_slice_proxy22[31:24]};
assign soc_videooverlaysoc_core_arp_depacketizer_source_param_sender_mac = {vns_slice_proxy31[7:0], vns_slice_proxy30[15:8], vns_slice_proxy29[23:16], vns_slice_proxy28[31:24], vns_slice_proxy27[39:32], vns_slice_proxy26[47:40]};
assign soc_videooverlaysoc_core_arp_depacketizer_source_param_target_ip = {vns_slice_proxy35[7:0], vns_slice_proxy34[15:8], vns_slice_proxy33[23:16], vns_slice_proxy32[31:24]};
assign soc_videooverlaysoc_core_arp_depacketizer_source_param_target_mac = {vns_slice_proxy41[7:0], vns_slice_proxy40[15:8], vns_slice_proxy39[23:16], vns_slice_proxy38[31:24], vns_slice_proxy37[39:32], vns_slice_proxy36[47:40]};
always @(*) begin
	soc_videooverlaysoc_core_arp_depacketizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_arp_depacketizer_counter_ce <= 1'd0;
	soc_videooverlaysoc_core_arp_depacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_arp_depacketizer_source_valid <= 1'd0;
	vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_next_state <= 2'd0;
	soc_videooverlaysoc_core_arp_depacketizer_shift <= 1'd0;
	vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_next_state <= vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_state;
	case (vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_core_arp_depacketizer_sink_ready <= 1'd1;
			if (soc_videooverlaysoc_core_arp_depacketizer_sink_valid) begin
				soc_videooverlaysoc_core_arp_depacketizer_counter_ce <= 1'd1;
				soc_videooverlaysoc_core_arp_depacketizer_shift <= 1'd1;
				if ((soc_videooverlaysoc_core_arp_depacketizer_counter == 5'd26)) begin
					vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_arp_depacketizer_sink_ready <= soc_videooverlaysoc_core_arp_depacketizer_source_ready;
			soc_videooverlaysoc_core_arp_depacketizer_source_valid <= (soc_videooverlaysoc_core_arp_depacketizer_sink_valid | soc_videooverlaysoc_core_arp_depacketizer_no_payload);
			if (((soc_videooverlaysoc_core_arp_depacketizer_source_valid & soc_videooverlaysoc_core_arp_depacketizer_source_ready) & soc_videooverlaysoc_core_arp_depacketizer_source_last)) begin
				vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_arp_depacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_arp_depacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_arp_depacketizer_sink_valid) begin
				soc_videooverlaysoc_core_arp_depacketizer_shift <= 1'd1;
				vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_arp_depacketizer_is_el = ((~(vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_state == 2'd2)) & (vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_next_state == 2'd2));
always @(*) begin
	soc_videooverlaysoc_core_arp_source_source_payload_reply <= 1'd0;
	soc_videooverlaysoc_core_arp_source_source_payload_request <= 1'd0;
	vns_clockdomainsrenamer1_liteetharprx_fsm_next_state <= 2'd0;
	soc_videooverlaysoc_core_arp_source_source_valid <= 1'd0;
	soc_videooverlaysoc_core_arp_depacketizer_source_ready <= 1'd0;
	vns_clockdomainsrenamer1_liteetharprx_fsm_next_state <= vns_clockdomainsrenamer1_liteetharprx_fsm_state;
	case (vns_clockdomainsrenamer1_liteetharprx_fsm_state)
		1'd1: begin
			if (soc_videooverlaysoc_core_arp_valid) begin
				soc_videooverlaysoc_core_arp_source_source_valid <= 1'd1;
				soc_videooverlaysoc_core_arp_source_source_payload_reply <= soc_videooverlaysoc_core_arp_reply;
				soc_videooverlaysoc_core_arp_source_source_payload_request <= soc_videooverlaysoc_core_arp_request;
			end
			vns_clockdomainsrenamer1_liteetharprx_fsm_next_state <= 2'd2;
		end
		2'd2: begin
			soc_videooverlaysoc_core_arp_depacketizer_source_ready <= 1'd1;
			if ((soc_videooverlaysoc_core_arp_depacketizer_source_valid & soc_videooverlaysoc_core_arp_depacketizer_source_last)) begin
				vns_clockdomainsrenamer1_liteetharprx_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_arp_depacketizer_source_ready <= 1'd1;
			if (soc_videooverlaysoc_core_arp_depacketizer_source_valid) begin
				soc_videooverlaysoc_core_arp_depacketizer_source_ready <= 1'd0;
				vns_clockdomainsrenamer1_liteetharprx_fsm_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_arp_table_request_timer_wait = (soc_videooverlaysoc_core_arp_table_request_pending & (~soc_videooverlaysoc_core_arp_table_request_counter_ce));
assign soc_videooverlaysoc_core_arp_table_cached_timer_wait = (~soc_videooverlaysoc_core_arp_table_update);
assign soc_videooverlaysoc_core_arp_table_response_payload_mac_address = soc_videooverlaysoc_core_arp_table_cached_mac_address;
assign soc_videooverlaysoc_core_arp_table_request_timer_done = (soc_videooverlaysoc_core_arp_table_request_timer_count == 1'd0);
assign soc_videooverlaysoc_core_arp_table_cached_timer_done = (soc_videooverlaysoc_core_arp_table_cached_timer_count == 1'd0);
always @(*) begin
	soc_videooverlaysoc_core_arp_table_source_payload_reply <= 1'd0;
	soc_videooverlaysoc_core_arp_table_request_pending_clr <= 1'd0;
	soc_videooverlaysoc_core_arp_table_source_payload_request <= 1'd0;
	soc_videooverlaysoc_core_arp_table_update <= 1'd0;
	soc_videooverlaysoc_core_arp_table_source_payload_ip_address <= 32'd0;
	soc_videooverlaysoc_core_arp_table_request_pending_set <= 1'd0;
	soc_videooverlaysoc_core_arp_table_source_payload_mac_address <= 48'd0;
	soc_videooverlaysoc_core_arp_table_response_payload_failed <= 1'd0;
	soc_videooverlaysoc_core_arp_table_request_ip_address_reset <= 1'd0;
	soc_videooverlaysoc_core_arp_table_request_ready <= 1'd0;
	soc_videooverlaysoc_core_arp_table_request_ip_address_update <= 1'd0;
	vns_clockdomainsrenamer1_next_state1 <= 3'd0;
	soc_videooverlaysoc_core_arp_table_response_valid <= 1'd0;
	soc_videooverlaysoc_core_arp_table_source_valid <= 1'd0;
	soc_videooverlaysoc_core_arp_table_request_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_arp_table_request_counter_ce <= 1'd0;
	if ((soc_videooverlaysoc_core_arp_table_request_counter == 3'd7)) begin
		soc_videooverlaysoc_core_arp_table_response_payload_failed <= 1'd1;
		soc_videooverlaysoc_core_arp_table_request_counter_reset <= 1'd1;
		soc_videooverlaysoc_core_arp_table_request_pending_clr <= 1'd1;
	end
	vns_clockdomainsrenamer1_next_state1 <= vns_clockdomainsrenamer1_state1;
	case (vns_clockdomainsrenamer1_state1)
		1'd1: begin
			soc_videooverlaysoc_core_arp_table_source_valid <= 1'd1;
			soc_videooverlaysoc_core_arp_table_source_payload_reply <= 1'd1;
			soc_videooverlaysoc_core_arp_table_source_payload_ip_address <= soc_videooverlaysoc_core_arp_table_sink_payload_ip_address;
			soc_videooverlaysoc_core_arp_table_source_payload_mac_address <= soc_videooverlaysoc_core_arp_table_sink_payload_mac_address;
			if (soc_videooverlaysoc_core_arp_table_source_ready) begin
				vns_clockdomainsrenamer1_next_state1 <= 1'd0;
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_arp_table_request_pending_clr <= 1'd1;
			soc_videooverlaysoc_core_arp_table_update <= 1'd1;
			vns_clockdomainsrenamer1_next_state1 <= 2'd3;
		end
		2'd3: begin
			if (soc_videooverlaysoc_core_arp_table_cached_valid) begin
				if ((soc_videooverlaysoc_core_arp_table_request_ip_address == soc_videooverlaysoc_core_arp_table_cached_ip_address)) begin
					soc_videooverlaysoc_core_arp_table_request_ip_address_reset <= 1'd1;
					vns_clockdomainsrenamer1_next_state1 <= 3'd5;
				end else begin
					if ((soc_videooverlaysoc_core_arp_table_request_payload_ip_address == soc_videooverlaysoc_core_arp_table_cached_ip_address)) begin
						soc_videooverlaysoc_core_arp_table_request_ready <= soc_videooverlaysoc_core_arp_table_request_valid;
						vns_clockdomainsrenamer1_next_state1 <= 3'd5;
					end else begin
						soc_videooverlaysoc_core_arp_table_request_ip_address_update <= soc_videooverlaysoc_core_arp_table_request_valid;
						vns_clockdomainsrenamer1_next_state1 <= 3'd4;
					end
				end
			end else begin
				soc_videooverlaysoc_core_arp_table_request_ip_address_update <= soc_videooverlaysoc_core_arp_table_request_valid;
				vns_clockdomainsrenamer1_next_state1 <= 3'd4;
			end
		end
		3'd4: begin
			soc_videooverlaysoc_core_arp_table_source_valid <= 1'd1;
			soc_videooverlaysoc_core_arp_table_source_payload_request <= 1'd1;
			soc_videooverlaysoc_core_arp_table_source_payload_ip_address <= soc_videooverlaysoc_core_arp_table_request_ip_address;
			if (soc_videooverlaysoc_core_arp_table_source_ready) begin
				soc_videooverlaysoc_core_arp_table_request_counter_reset <= soc_videooverlaysoc_core_arp_table_request_valid;
				soc_videooverlaysoc_core_arp_table_request_counter_ce <= 1'd1;
				soc_videooverlaysoc_core_arp_table_request_pending_set <= 1'd1;
				soc_videooverlaysoc_core_arp_table_request_ready <= 1'd1;
				vns_clockdomainsrenamer1_next_state1 <= 1'd0;
			end
		end
		3'd5: begin
			soc_videooverlaysoc_core_arp_table_response_valid <= 1'd1;
			if (soc_videooverlaysoc_core_arp_table_response_ready) begin
				vns_clockdomainsrenamer1_next_state1 <= 1'd0;
			end
		end
		default: begin
			if ((soc_videooverlaysoc_core_arp_table_sink_valid & soc_videooverlaysoc_core_arp_table_sink_payload_request)) begin
				vns_clockdomainsrenamer1_next_state1 <= 1'd1;
			end else begin
				if (((soc_videooverlaysoc_core_arp_table_sink_valid & soc_videooverlaysoc_core_arp_table_sink_payload_reply) & soc_videooverlaysoc_core_arp_table_request_pending)) begin
					vns_clockdomainsrenamer1_next_state1 <= 2'd2;
				end else begin
					if ((soc_videooverlaysoc_core_arp_table_request_counter == 3'd7)) begin
						vns_clockdomainsrenamer1_next_state1 <= 3'd5;
					end else begin
						if ((soc_videooverlaysoc_core_arp_table_request_valid | (soc_videooverlaysoc_core_arp_table_request_pending & soc_videooverlaysoc_core_arp_table_request_timer_done))) begin
							vns_clockdomainsrenamer1_next_state1 <= 2'd3;
						end
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_ip_mac_port_sink_valid = soc_videooverlaysoc_core_ip_tx_source_valid;
assign soc_videooverlaysoc_core_ip_tx_source_ready = soc_videooverlaysoc_core_ip_mac_port_sink_ready;
assign soc_videooverlaysoc_core_ip_mac_port_sink_first = soc_videooverlaysoc_core_ip_tx_source_first;
assign soc_videooverlaysoc_core_ip_mac_port_sink_last = soc_videooverlaysoc_core_ip_tx_source_last;
assign soc_videooverlaysoc_core_ip_mac_port_sink_payload_ethernet_type = soc_videooverlaysoc_core_ip_tx_source_payload_ethernet_type;
assign soc_videooverlaysoc_core_ip_mac_port_sink_payload_sender_mac = soc_videooverlaysoc_core_ip_tx_source_payload_sender_mac;
assign soc_videooverlaysoc_core_ip_mac_port_sink_payload_target_mac = soc_videooverlaysoc_core_ip_tx_source_payload_target_mac;
assign soc_videooverlaysoc_core_ip_mac_port_sink_payload_data = soc_videooverlaysoc_core_ip_tx_source_payload_data;
assign soc_videooverlaysoc_core_ip_mac_port_sink_payload_last_be = soc_videooverlaysoc_core_ip_tx_source_payload_last_be;
assign soc_videooverlaysoc_core_ip_mac_port_sink_payload_error = soc_videooverlaysoc_core_ip_tx_source_payload_error;
assign soc_videooverlaysoc_core_ip_rx_sink_sink_valid = soc_videooverlaysoc_core_ip_mac_port_source_valid;
assign soc_videooverlaysoc_core_ip_mac_port_source_ready = soc_videooverlaysoc_core_ip_rx_sink_sink_ready;
assign soc_videooverlaysoc_core_ip_rx_sink_sink_first = soc_videooverlaysoc_core_ip_mac_port_source_first;
assign soc_videooverlaysoc_core_ip_rx_sink_sink_last = soc_videooverlaysoc_core_ip_mac_port_source_last;
assign soc_videooverlaysoc_core_ip_rx_sink_sink_payload_ethernet_type = soc_videooverlaysoc_core_ip_mac_port_source_payload_ethernet_type;
assign soc_videooverlaysoc_core_ip_rx_sink_sink_payload_sender_mac = soc_videooverlaysoc_core_ip_mac_port_source_payload_sender_mac;
assign soc_videooverlaysoc_core_ip_rx_sink_sink_payload_target_mac = soc_videooverlaysoc_core_ip_mac_port_source_payload_target_mac;
assign soc_videooverlaysoc_core_ip_rx_sink_sink_payload_data = soc_videooverlaysoc_core_ip_mac_port_source_payload_data;
assign soc_videooverlaysoc_core_ip_rx_sink_sink_payload_last_be = soc_videooverlaysoc_core_ip_mac_port_source_payload_last_be;
assign soc_videooverlaysoc_core_ip_rx_sink_sink_payload_error = soc_videooverlaysoc_core_ip_mac_port_source_payload_error;
assign soc_videooverlaysoc_core_ip_tx_sink_valid = soc_videooverlaysoc_core_ip_crossbar_source_valid;
assign soc_videooverlaysoc_core_ip_crossbar_source_ready = soc_videooverlaysoc_core_ip_tx_sink_ready;
assign soc_videooverlaysoc_core_ip_tx_sink_first = soc_videooverlaysoc_core_ip_crossbar_source_first;
assign soc_videooverlaysoc_core_ip_tx_sink_last = soc_videooverlaysoc_core_ip_crossbar_source_last;
assign soc_videooverlaysoc_core_ip_tx_sink_payload_data = soc_videooverlaysoc_core_ip_crossbar_source_payload_data;
assign soc_videooverlaysoc_core_ip_tx_sink_payload_error = soc_videooverlaysoc_core_ip_crossbar_source_payload_error;
assign soc_videooverlaysoc_core_ip_tx_sink_param_length = soc_videooverlaysoc_core_ip_crossbar_source_param_length;
assign soc_videooverlaysoc_core_ip_tx_sink_param_protocol = soc_videooverlaysoc_core_ip_crossbar_source_param_protocol;
assign soc_videooverlaysoc_core_ip_tx_sink_param_ip_address = soc_videooverlaysoc_core_ip_crossbar_source_param_ip_address;
assign soc_videooverlaysoc_core_ip_crossbar_sink_valid = soc_videooverlaysoc_core_ip_rx_source_source_valid;
assign soc_videooverlaysoc_core_ip_rx_source_source_ready = soc_videooverlaysoc_core_ip_crossbar_sink_ready;
assign soc_videooverlaysoc_core_ip_crossbar_sink_first = soc_videooverlaysoc_core_ip_rx_source_source_first;
assign soc_videooverlaysoc_core_ip_crossbar_sink_last = soc_videooverlaysoc_core_ip_rx_source_source_last;
assign soc_videooverlaysoc_core_ip_crossbar_sink_payload_data = soc_videooverlaysoc_core_ip_rx_source_source_payload_data;
assign soc_videooverlaysoc_core_ip_crossbar_sink_payload_error = soc_videooverlaysoc_core_ip_rx_source_source_payload_error;
assign soc_videooverlaysoc_core_ip_crossbar_sink_param_length = soc_videooverlaysoc_core_ip_rx_source_source_param_length;
assign soc_videooverlaysoc_core_ip_crossbar_sink_param_protocol = soc_videooverlaysoc_core_ip_rx_source_source_param_protocol;
assign soc_videooverlaysoc_core_ip_crossbar_sink_param_ip_address = soc_videooverlaysoc_core_ip_rx_source_source_param_ip_address;
assign soc_videooverlaysoc_core_ip_tx_ce = soc_videooverlaysoc_core_ip_tx_sink_valid;
assign soc_videooverlaysoc_core_ip_tx_reset = ((soc_videooverlaysoc_core_ip_tx_source_valid & soc_videooverlaysoc_core_ip_tx_source_last) & soc_videooverlaysoc_core_ip_tx_source_ready);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_valid = (soc_videooverlaysoc_core_ip_tx_sink_valid & soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_last = soc_videooverlaysoc_core_ip_tx_sink_last;
assign soc_videooverlaysoc_core_ip_tx_sink_ready = (soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_ready & soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_target_ip = soc_videooverlaysoc_core_ip_tx_sink_param_ip_address;
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_protocol = soc_videooverlaysoc_core_ip_tx_sink_param_protocol;
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_total_length = (soc_videooverlaysoc_core_ip_tx_sink_param_length + 5'd20);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_version = 3'd4;
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_ihl = 3'd5;
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_identification = 1'd0;
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_ttl = 8'd128;
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_sender_ip = 28'd167774978;
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_payload_data = soc_videooverlaysoc_core_ip_tx_sink_payload_data;
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header = soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header;
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_checksum = soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_value;
assign soc_videooverlaysoc_core_arp_table_request_payload_ip_address = soc_videooverlaysoc_core_ip_tx_sink_param_ip_address;
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next0 = (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header[15:0]);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next1 = (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next0 + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header[31:16]);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next2 = (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next1 + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header[47:32]);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next3 = (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next2 + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header[63:48]);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next4 = (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next3 + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header[79:64]);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next5 = (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next4 + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header[111:96]);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next6 = (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next5 + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header[127:112]);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next7 = (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next6 + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header[143:128]);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next8 = (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next7 + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_header[159:144]);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_value = (~{soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next8[7:0], soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next8[15:8]});
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_counter_ce = (~soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done);
assign soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done = (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_counter == 4'd9);
always @(*) begin
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header <= 160'd0;
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header[95:80] <= {soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_checksum[7:0], soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_checksum[15:8]};
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header[47:32] <= {soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_identification[7:0], soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_identification[15:8]};
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header[3:0] <= {soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_ihl[3:0]};
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header[79:72] <= {soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_protocol[7:0]};
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header[127:96] <= {soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_sender_ip[7:0], soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_sender_ip[15:8], soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_sender_ip[23:16], soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_sender_ip[31:24]};
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header[159:128] <= {soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_target_ip[7:0], soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_target_ip[15:8], soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_target_ip[23:16], soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_target_ip[31:24]};
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header[31:16] <= {soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_total_length[7:0], soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_total_length[15:8]};
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header[71:64] <= {soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_ttl[7:0]};
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header[7:4] <= {soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_param_version[3:0]};
end
assign soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_error = soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_payload_error;
always @(*) begin
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_load <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_shift <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter_ce <= 1'd0;
	vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_next_state <= 2'd0;
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_last <= 1'd0;
	vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_next_state <= vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_state;
	case (vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_state)
		1'd1: begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid <= 1'd1;
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_last <= 1'd0;
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_data <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header_reg[15:8];
			if ((soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid & soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_ready)) begin
				soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_shift <= 1'd1;
				soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter_ce <= 1'd1;
				if ((soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter == 5'd18)) begin
					vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_valid;
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_last <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_last;
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_data <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_payload_data;
			if ((soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid & soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_ready)) begin
				soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_ready <= 1'd1;
				if (soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_last) begin
					vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_valid) begin
				soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_sink_ready <= 1'd0;
				soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid <= 1'd1;
				soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_last <= 1'd0;
				soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_data <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header[7:0];
				if ((soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid & soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_ready)) begin
					soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_load <= 1'd1;
					vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_next_state <= 1'd1;
				end
			end
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_core_ip_tx_target_unreachable <= 1'd0;
	vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_next_state <= 3'd0;
	soc_videooverlaysoc_core_arp_table_request_valid <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_source_valid <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_source_first <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_source_last <= 1'd0;
	soc_videooverlaysoc_core_arp_table_response_ready <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_ready <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_source_payload_ethernet_type <= 16'd0;
	soc_videooverlaysoc_core_ip_tx_source_payload_sender_mac <= 48'd0;
	soc_videooverlaysoc_core_ip_tx_source_payload_target_mac <= 48'd0;
	soc_videooverlaysoc_core_ip_tx_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_ip_tx_source_payload_last_be <= 1'd0;
	soc_videooverlaysoc_core_ip_tx_source_payload_error <= 1'd0;
	vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_next_state <= vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_state;
	case (vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_state)
		1'd1: begin
			soc_videooverlaysoc_core_arp_table_request_valid <= 1'd1;
			if ((soc_videooverlaysoc_core_arp_table_request_valid & soc_videooverlaysoc_core_arp_table_request_ready)) begin
				vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (soc_videooverlaysoc_core_arp_table_response_valid) begin
				soc_videooverlaysoc_core_arp_table_response_ready <= 1'd1;
				if (soc_videooverlaysoc_core_arp_table_response_payload_failed) begin
					soc_videooverlaysoc_core_ip_tx_target_unreachable <= 1'd1;
					vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_next_state <= 3'd4;
				end else begin
					vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_next_state <= 2'd3;
				end
			end
		end
		2'd3: begin
			soc_videooverlaysoc_core_ip_tx_source_valid <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid;
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_ready <= soc_videooverlaysoc_core_ip_tx_source_ready;
			soc_videooverlaysoc_core_ip_tx_source_first <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_first;
			soc_videooverlaysoc_core_ip_tx_source_last <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_last;
			soc_videooverlaysoc_core_ip_tx_source_payload_ethernet_type <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_ethernet_type;
			soc_videooverlaysoc_core_ip_tx_source_payload_sender_mac <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_sender_mac;
			soc_videooverlaysoc_core_ip_tx_source_payload_target_mac <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_target_mac;
			soc_videooverlaysoc_core_ip_tx_source_payload_data <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_data;
			soc_videooverlaysoc_core_ip_tx_source_payload_last_be <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_last_be;
			soc_videooverlaysoc_core_ip_tx_source_payload_error <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_payload_error;
			soc_videooverlaysoc_core_ip_tx_source_payload_ethernet_type <= 12'd2048;
			soc_videooverlaysoc_core_ip_tx_source_payload_target_mac <= soc_videooverlaysoc_core_ip_tx_target_mac;
			soc_videooverlaysoc_core_ip_tx_source_payload_sender_mac <= 45'd21127783889598;
			if (((soc_videooverlaysoc_core_ip_tx_source_valid & soc_videooverlaysoc_core_ip_tx_source_last) & soc_videooverlaysoc_core_ip_tx_source_ready)) begin
				vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_next_state <= 1'd0;
			end
		end
		3'd4: begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_ready <= 1'd1;
			if (((soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid & soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_last) & soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_ready)) begin
				vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_ready <= 1'd1;
			if (soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_valid) begin
				soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_source_ready <= 1'd0;
				vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_ip_rx_depacketizer_sink_valid = soc_videooverlaysoc_core_ip_rx_sink_sink_valid;
assign soc_videooverlaysoc_core_ip_rx_sink_sink_ready = soc_videooverlaysoc_core_ip_rx_depacketizer_sink_ready;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_sink_first = soc_videooverlaysoc_core_ip_rx_sink_sink_first;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_sink_last = soc_videooverlaysoc_core_ip_rx_sink_sink_last;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_ethernet_type = soc_videooverlaysoc_core_ip_rx_sink_sink_payload_ethernet_type;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_sender_mac = soc_videooverlaysoc_core_ip_rx_sink_sink_payload_sender_mac;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_target_mac = soc_videooverlaysoc_core_ip_rx_sink_sink_payload_target_mac;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_data = soc_videooverlaysoc_core_ip_rx_sink_sink_payload_data;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_last_be = soc_videooverlaysoc_core_ip_rx_sink_sink_payload_last_be;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_error = soc_videooverlaysoc_core_ip_rx_sink_sink_payload_error;
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header = soc_videooverlaysoc_core_ip_rx_depacketizer_header;
assign soc_videooverlaysoc_core_ip_rx_reset = (~soc_videooverlaysoc_core_ip_rx_depacketizer_source_valid);
assign soc_videooverlaysoc_core_ip_rx_ce = 1'd1;
assign soc_videooverlaysoc_core_ip_rx_source_source_last = soc_videooverlaysoc_core_ip_rx_depacketizer_source_last;
assign soc_videooverlaysoc_core_ip_rx_source_source_param_length = (soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_total_length - 5'd20);
assign soc_videooverlaysoc_core_ip_rx_source_source_param_protocol = soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_protocol;
assign soc_videooverlaysoc_core_ip_rx_source_source_param_ip_address = soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_sender_ip;
assign soc_videooverlaysoc_core_ip_rx_source_source_payload_data = soc_videooverlaysoc_core_ip_rx_depacketizer_source_payload_data;
assign soc_videooverlaysoc_core_ip_rx_source_source_payload_error = soc_videooverlaysoc_core_ip_rx_depacketizer_source_payload_error;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_header = soc_videooverlaysoc_core_ip_rx_depacketizer_header_reg;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_payload_error = soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_error;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_last = (soc_videooverlaysoc_core_ip_rx_depacketizer_sink_last | soc_videooverlaysoc_core_ip_rx_depacketizer_no_payload);
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_payload_data = soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_data;
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_checksum = {vns_slice_proxy43[7:0], vns_slice_proxy42[15:8]};
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_identification = {vns_slice_proxy45[7:0], vns_slice_proxy44[15:8]};
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_ihl = {vns_slice_proxy46[3:0]};
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_protocol = {vns_slice_proxy47[7:0]};
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_sender_ip = {vns_slice_proxy51[7:0], vns_slice_proxy50[15:8], vns_slice_proxy49[23:16], vns_slice_proxy48[31:24]};
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_target_ip = {vns_slice_proxy55[7:0], vns_slice_proxy54[15:8], vns_slice_proxy53[23:16], vns_slice_proxy52[31:24]};
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_total_length = {vns_slice_proxy57[7:0], vns_slice_proxy56[15:8]};
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_ttl = {vns_slice_proxy58[7:0]};
assign soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_version = {vns_slice_proxy59[3:0]};
always @(*) begin
	soc_videooverlaysoc_core_ip_rx_depacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_ip_rx_depacketizer_source_valid <= 1'd0;
	soc_videooverlaysoc_core_ip_rx_depacketizer_shift <= 1'd0;
	soc_videooverlaysoc_core_ip_rx_depacketizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_ip_rx_depacketizer_counter_ce <= 1'd0;
	vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_next_state <= 2'd0;
	vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_next_state <= vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_state;
	case (vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_core_ip_rx_depacketizer_sink_ready <= 1'd1;
			if (soc_videooverlaysoc_core_ip_rx_depacketizer_sink_valid) begin
				soc_videooverlaysoc_core_ip_rx_depacketizer_counter_ce <= 1'd1;
				soc_videooverlaysoc_core_ip_rx_depacketizer_shift <= 1'd1;
				if ((soc_videooverlaysoc_core_ip_rx_depacketizer_counter == 5'd18)) begin
					vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_ip_rx_depacketizer_sink_ready <= soc_videooverlaysoc_core_ip_rx_depacketizer_source_ready;
			soc_videooverlaysoc_core_ip_rx_depacketizer_source_valid <= (soc_videooverlaysoc_core_ip_rx_depacketizer_sink_valid | soc_videooverlaysoc_core_ip_rx_depacketizer_no_payload);
			if (((soc_videooverlaysoc_core_ip_rx_depacketizer_source_valid & soc_videooverlaysoc_core_ip_rx_depacketizer_source_ready) & soc_videooverlaysoc_core_ip_rx_depacketizer_source_last)) begin
				vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_ip_rx_depacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_ip_rx_depacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_ip_rx_depacketizer_sink_valid) begin
				soc_videooverlaysoc_core_ip_rx_depacketizer_shift <= 1'd1;
				vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_ip_rx_depacketizer_is_el = ((~(vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_state == 2'd2)) & (vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_next_state == 2'd2));
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next0 = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header[15:0]);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next1 = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next0 + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header[31:16]);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next2 = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next1 + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header[47:32]);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next3 = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next2 + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header[63:48]);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next4 = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next3 + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header[79:64]);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next5 = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next4 + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header[95:80]);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next6 = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next5 + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header[111:96]);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next7 = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next6 + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header[127:112]);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next8 = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next7 + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header[143:128]);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next9 = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next8 + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_header[159:144]);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_value = (~{soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next9[7:0], soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next9[15:8]});
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_counter_ce = (~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done);
assign soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done = (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_counter == 4'd11);
always @(*) begin
	soc_videooverlaysoc_core_ip_rx_depacketizer_source_ready <= 1'd0;
	vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_next_state <= 2'd0;
	soc_videooverlaysoc_core_ip_rx_source_source_valid <= 1'd0;
	vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_next_state <= vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_state;
	case (vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_state)
		1'd1: begin
			if (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done) begin
				if (soc_videooverlaysoc_core_ip_rx_valid) begin
					vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_next_state <= 2'd2;
				end else begin
					vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_ip_rx_source_source_valid <= soc_videooverlaysoc_core_ip_rx_depacketizer_source_valid;
			soc_videooverlaysoc_core_ip_rx_depacketizer_source_ready <= soc_videooverlaysoc_core_ip_rx_source_source_ready;
			if (((soc_videooverlaysoc_core_ip_rx_source_source_valid & soc_videooverlaysoc_core_ip_rx_source_source_last) & soc_videooverlaysoc_core_ip_rx_source_source_ready)) begin
				vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_next_state <= 1'd0;
			end
		end
		2'd3: begin
			soc_videooverlaysoc_core_ip_rx_depacketizer_source_ready <= 1'd1;
			if (((soc_videooverlaysoc_core_ip_rx_depacketizer_source_valid & soc_videooverlaysoc_core_ip_rx_depacketizer_source_last) & soc_videooverlaysoc_core_ip_rx_depacketizer_source_ready)) begin
				vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_ip_rx_depacketizer_source_ready <= 1'd1;
			if (soc_videooverlaysoc_core_ip_rx_depacketizer_source_valid) begin
				soc_videooverlaysoc_core_ip_rx_depacketizer_source_ready <= 1'd0;
				vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_next_state <= 1'd1;
			end
		end
	endcase
end
always @(*) begin
	vns_clockdomainsrenamer1_liteethip_sel0 <= 2'd0;
	case (soc_videooverlaysoc_core_ip_crossbar_sink_param_protocol)
		1'd1: begin
			vns_clockdomainsrenamer1_liteethip_sel0 <= 1'd1;
		end
		5'd17: begin
			vns_clockdomainsrenamer1_liteethip_sel0 <= 2'd2;
		end
		default: begin
			vns_clockdomainsrenamer1_liteethip_sel0 <= 1'd0;
		end
	endcase
end
always @(*) begin
	vns_clockdomainsrenamer1_liteethip_request <= 2'd0;
	vns_clockdomainsrenamer1_liteethip_request[0] <= vns_clockdomainsrenamer1_liteethip_status0_ongoing0;
	vns_clockdomainsrenamer1_liteethip_request[1] <= vns_clockdomainsrenamer1_liteethip_status1_ongoing0;
end
always @(*) begin
	soc_videooverlaysoc_core_ip_crossbar_source_valid <= 1'd0;
	soc_videooverlaysoc_core_ip_port_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_ip_crossbar_source_first <= 1'd0;
	soc_videooverlaysoc_core_ip_crossbar_source_last <= 1'd0;
	soc_videooverlaysoc_core_icmp_ip_port_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_ip_crossbar_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_ip_crossbar_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_ip_crossbar_source_param_length <= 16'd0;
	soc_videooverlaysoc_core_ip_crossbar_source_param_protocol <= 8'd0;
	soc_videooverlaysoc_core_ip_crossbar_source_param_ip_address <= 32'd0;
	case (vns_clockdomainsrenamer1_liteethip_grant)
		1'd0: begin
			soc_videooverlaysoc_core_ip_crossbar_source_valid <= soc_videooverlaysoc_core_icmp_ip_port_sink_valid;
			soc_videooverlaysoc_core_icmp_ip_port_sink_ready <= soc_videooverlaysoc_core_ip_crossbar_source_ready;
			soc_videooverlaysoc_core_ip_crossbar_source_first <= soc_videooverlaysoc_core_icmp_ip_port_sink_first;
			soc_videooverlaysoc_core_ip_crossbar_source_last <= soc_videooverlaysoc_core_icmp_ip_port_sink_last;
			soc_videooverlaysoc_core_ip_crossbar_source_payload_data <= soc_videooverlaysoc_core_icmp_ip_port_sink_payload_data;
			soc_videooverlaysoc_core_ip_crossbar_source_payload_error <= soc_videooverlaysoc_core_icmp_ip_port_sink_payload_error;
			soc_videooverlaysoc_core_ip_crossbar_source_param_length <= soc_videooverlaysoc_core_icmp_ip_port_sink_param_length;
			soc_videooverlaysoc_core_ip_crossbar_source_param_protocol <= soc_videooverlaysoc_core_icmp_ip_port_sink_param_protocol;
			soc_videooverlaysoc_core_ip_crossbar_source_param_ip_address <= soc_videooverlaysoc_core_icmp_ip_port_sink_param_ip_address;
		end
		1'd1: begin
			soc_videooverlaysoc_core_ip_crossbar_source_valid <= soc_videooverlaysoc_core_ip_port_sink_valid;
			soc_videooverlaysoc_core_ip_port_sink_ready <= soc_videooverlaysoc_core_ip_crossbar_source_ready;
			soc_videooverlaysoc_core_ip_crossbar_source_first <= soc_videooverlaysoc_core_ip_port_sink_first;
			soc_videooverlaysoc_core_ip_crossbar_source_last <= soc_videooverlaysoc_core_ip_port_sink_last;
			soc_videooverlaysoc_core_ip_crossbar_source_payload_data <= soc_videooverlaysoc_core_ip_port_sink_payload_data;
			soc_videooverlaysoc_core_ip_crossbar_source_payload_error <= soc_videooverlaysoc_core_ip_port_sink_payload_error;
			soc_videooverlaysoc_core_ip_crossbar_source_param_length <= soc_videooverlaysoc_core_ip_port_sink_param_length;
			soc_videooverlaysoc_core_ip_crossbar_source_param_protocol <= soc_videooverlaysoc_core_ip_port_sink_param_protocol;
			soc_videooverlaysoc_core_ip_crossbar_source_param_ip_address <= soc_videooverlaysoc_core_ip_port_sink_param_ip_address;
		end
	endcase
end
always @(*) begin
	vns_clockdomainsrenamer1_liteethip_status0_last <= 1'd0;
	if (soc_videooverlaysoc_core_icmp_ip_port_sink_valid) begin
		vns_clockdomainsrenamer1_liteethip_status0_last <= (soc_videooverlaysoc_core_icmp_ip_port_sink_last & soc_videooverlaysoc_core_icmp_ip_port_sink_ready);
	end
end
assign vns_clockdomainsrenamer1_liteethip_status0_ongoing0 = ((soc_videooverlaysoc_core_icmp_ip_port_sink_valid | vns_clockdomainsrenamer1_liteethip_status0_ongoing1) & (~vns_clockdomainsrenamer1_liteethip_status0_last));
always @(*) begin
	vns_clockdomainsrenamer1_liteethip_status1_last <= 1'd0;
	if (soc_videooverlaysoc_core_ip_port_sink_valid) begin
		vns_clockdomainsrenamer1_liteethip_status1_last <= (soc_videooverlaysoc_core_ip_port_sink_last & soc_videooverlaysoc_core_ip_port_sink_ready);
	end
end
assign vns_clockdomainsrenamer1_liteethip_status1_ongoing0 = ((soc_videooverlaysoc_core_ip_port_sink_valid | vns_clockdomainsrenamer1_liteethip_status1_ongoing1) & (~vns_clockdomainsrenamer1_liteethip_status1_last));
always @(*) begin
	vns_clockdomainsrenamer1_liteethip_sel1 <= 2'd0;
	if (vns_clockdomainsrenamer1_liteethip_first) begin
		vns_clockdomainsrenamer1_liteethip_sel1 <= vns_clockdomainsrenamer1_liteethip_sel0;
	end else begin
		vns_clockdomainsrenamer1_liteethip_sel1 <= vns_clockdomainsrenamer1_liteethip_sel_ongoing;
	end
end
always @(*) begin
	soc_videooverlaysoc_core_ip_port_source_valid <= 1'd0;
	soc_videooverlaysoc_core_ip_port_source_first <= 1'd0;
	soc_videooverlaysoc_core_icmp_ip_port_source_valid <= 1'd0;
	soc_videooverlaysoc_core_ip_port_source_last <= 1'd0;
	soc_videooverlaysoc_core_ip_port_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_ip_port_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_icmp_ip_port_source_first <= 1'd0;
	soc_videooverlaysoc_core_icmp_ip_port_source_last <= 1'd0;
	soc_videooverlaysoc_core_ip_port_source_param_length <= 16'd0;
	soc_videooverlaysoc_core_icmp_ip_port_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_ip_port_source_param_protocol <= 8'd0;
	soc_videooverlaysoc_core_icmp_ip_port_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_ip_port_source_param_ip_address <= 32'd0;
	soc_videooverlaysoc_core_icmp_ip_port_source_param_length <= 16'd0;
	soc_videooverlaysoc_core_icmp_ip_port_source_param_protocol <= 8'd0;
	soc_videooverlaysoc_core_icmp_ip_port_source_param_ip_address <= 32'd0;
	soc_videooverlaysoc_core_ip_crossbar_sink_ready <= 1'd0;
	case (vns_clockdomainsrenamer1_liteethip_sel1)
		1'd1: begin
			soc_videooverlaysoc_core_icmp_ip_port_source_valid <= soc_videooverlaysoc_core_ip_crossbar_sink_valid;
			soc_videooverlaysoc_core_ip_crossbar_sink_ready <= soc_videooverlaysoc_core_icmp_ip_port_source_ready;
			soc_videooverlaysoc_core_icmp_ip_port_source_first <= soc_videooverlaysoc_core_ip_crossbar_sink_first;
			soc_videooverlaysoc_core_icmp_ip_port_source_last <= soc_videooverlaysoc_core_ip_crossbar_sink_last;
			soc_videooverlaysoc_core_icmp_ip_port_source_payload_data <= soc_videooverlaysoc_core_ip_crossbar_sink_payload_data;
			soc_videooverlaysoc_core_icmp_ip_port_source_payload_error <= soc_videooverlaysoc_core_ip_crossbar_sink_payload_error;
			soc_videooverlaysoc_core_icmp_ip_port_source_param_length <= soc_videooverlaysoc_core_ip_crossbar_sink_param_length;
			soc_videooverlaysoc_core_icmp_ip_port_source_param_protocol <= soc_videooverlaysoc_core_ip_crossbar_sink_param_protocol;
			soc_videooverlaysoc_core_icmp_ip_port_source_param_ip_address <= soc_videooverlaysoc_core_ip_crossbar_sink_param_ip_address;
		end
		2'd2: begin
			soc_videooverlaysoc_core_ip_port_source_valid <= soc_videooverlaysoc_core_ip_crossbar_sink_valid;
			soc_videooverlaysoc_core_ip_crossbar_sink_ready <= soc_videooverlaysoc_core_ip_port_source_ready;
			soc_videooverlaysoc_core_ip_port_source_first <= soc_videooverlaysoc_core_ip_crossbar_sink_first;
			soc_videooverlaysoc_core_ip_port_source_last <= soc_videooverlaysoc_core_ip_crossbar_sink_last;
			soc_videooverlaysoc_core_ip_port_source_payload_data <= soc_videooverlaysoc_core_ip_crossbar_sink_payload_data;
			soc_videooverlaysoc_core_ip_port_source_payload_error <= soc_videooverlaysoc_core_ip_crossbar_sink_payload_error;
			soc_videooverlaysoc_core_ip_port_source_param_length <= soc_videooverlaysoc_core_ip_crossbar_sink_param_length;
			soc_videooverlaysoc_core_ip_port_source_param_protocol <= soc_videooverlaysoc_core_ip_crossbar_sink_param_protocol;
			soc_videooverlaysoc_core_ip_port_source_param_ip_address <= soc_videooverlaysoc_core_ip_crossbar_sink_param_ip_address;
		end
		default: begin
			soc_videooverlaysoc_core_ip_crossbar_sink_ready <= 1'd1;
		end
	endcase
end
always @(*) begin
	vns_clockdomainsrenamer1_liteethip_last <= 1'd0;
	if (soc_videooverlaysoc_core_ip_crossbar_sink_valid) begin
		vns_clockdomainsrenamer1_liteethip_last <= (soc_videooverlaysoc_core_ip_crossbar_sink_last & soc_videooverlaysoc_core_ip_crossbar_sink_ready);
	end
end
assign vns_clockdomainsrenamer1_liteethip_ongoing0 = ((soc_videooverlaysoc_core_ip_crossbar_sink_valid | vns_clockdomainsrenamer1_liteethip_ongoing1) & (~vns_clockdomainsrenamer1_liteethip_last));
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_valid = soc_videooverlaysoc_core_icmp_rx_source_source_valid;
assign soc_videooverlaysoc_core_icmp_rx_source_source_ready = soc_videooverlaysoc_core_icmp_echo_sink_sink_ready;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_first = soc_videooverlaysoc_core_icmp_rx_source_source_first;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_last = soc_videooverlaysoc_core_icmp_rx_source_source_last;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_payload_data = soc_videooverlaysoc_core_icmp_rx_source_source_payload_data;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_payload_error = soc_videooverlaysoc_core_icmp_rx_source_source_payload_error;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_param_checksum = soc_videooverlaysoc_core_icmp_rx_source_source_param_checksum;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_param_code = soc_videooverlaysoc_core_icmp_rx_source_source_param_code;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_param_msgtype = soc_videooverlaysoc_core_icmp_rx_source_source_param_msgtype;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_param_quench = soc_videooverlaysoc_core_icmp_rx_source_source_param_quench;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_param_ip_address = soc_videooverlaysoc_core_icmp_rx_source_source_param_ip_address;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_param_length = soc_videooverlaysoc_core_icmp_rx_source_source_param_length;
assign soc_videooverlaysoc_core_icmp_tx_sink_valid = soc_videooverlaysoc_core_icmp_echo_source_source_valid;
assign soc_videooverlaysoc_core_icmp_echo_source_source_ready = soc_videooverlaysoc_core_icmp_tx_sink_ready;
assign soc_videooverlaysoc_core_icmp_tx_sink_first = soc_videooverlaysoc_core_icmp_echo_source_source_first;
assign soc_videooverlaysoc_core_icmp_tx_sink_last = soc_videooverlaysoc_core_icmp_echo_source_source_last;
assign soc_videooverlaysoc_core_icmp_tx_sink_payload_data = soc_videooverlaysoc_core_icmp_echo_source_source_payload_data;
assign soc_videooverlaysoc_core_icmp_tx_sink_payload_error = soc_videooverlaysoc_core_icmp_echo_source_source_payload_error;
assign soc_videooverlaysoc_core_icmp_tx_sink_param_checksum = soc_videooverlaysoc_core_icmp_echo_source_source_param_checksum;
assign soc_videooverlaysoc_core_icmp_tx_sink_param_code = soc_videooverlaysoc_core_icmp_echo_source_source_param_code;
assign soc_videooverlaysoc_core_icmp_tx_sink_param_msgtype = soc_videooverlaysoc_core_icmp_echo_source_source_param_msgtype;
assign soc_videooverlaysoc_core_icmp_tx_sink_param_quench = soc_videooverlaysoc_core_icmp_echo_source_source_param_quench;
assign soc_videooverlaysoc_core_icmp_tx_sink_param_ip_address = soc_videooverlaysoc_core_icmp_echo_source_source_param_ip_address;
assign soc_videooverlaysoc_core_icmp_tx_sink_param_length = soc_videooverlaysoc_core_icmp_echo_source_source_param_length;
assign soc_videooverlaysoc_core_icmp_ip_port_sink_valid = soc_videooverlaysoc_core_icmp_tx_source_valid;
assign soc_videooverlaysoc_core_icmp_tx_source_ready = soc_videooverlaysoc_core_icmp_ip_port_sink_ready;
assign soc_videooverlaysoc_core_icmp_ip_port_sink_first = soc_videooverlaysoc_core_icmp_tx_source_first;
assign soc_videooverlaysoc_core_icmp_ip_port_sink_last = soc_videooverlaysoc_core_icmp_tx_source_last;
assign soc_videooverlaysoc_core_icmp_ip_port_sink_payload_data = soc_videooverlaysoc_core_icmp_tx_source_payload_data;
assign soc_videooverlaysoc_core_icmp_ip_port_sink_payload_error = soc_videooverlaysoc_core_icmp_tx_source_payload_error;
assign soc_videooverlaysoc_core_icmp_ip_port_sink_param_length = soc_videooverlaysoc_core_icmp_tx_source_param_length;
assign soc_videooverlaysoc_core_icmp_ip_port_sink_param_protocol = soc_videooverlaysoc_core_icmp_tx_source_param_protocol;
assign soc_videooverlaysoc_core_icmp_ip_port_sink_param_ip_address = soc_videooverlaysoc_core_icmp_tx_source_param_ip_address;
assign soc_videooverlaysoc_core_icmp_rx_sink_sink_valid = soc_videooverlaysoc_core_icmp_ip_port_source_valid;
assign soc_videooverlaysoc_core_icmp_ip_port_source_ready = soc_videooverlaysoc_core_icmp_rx_sink_sink_ready;
assign soc_videooverlaysoc_core_icmp_rx_sink_sink_first = soc_videooverlaysoc_core_icmp_ip_port_source_first;
assign soc_videooverlaysoc_core_icmp_rx_sink_sink_last = soc_videooverlaysoc_core_icmp_ip_port_source_last;
assign soc_videooverlaysoc_core_icmp_rx_sink_sink_payload_data = soc_videooverlaysoc_core_icmp_ip_port_source_payload_data;
assign soc_videooverlaysoc_core_icmp_rx_sink_sink_payload_error = soc_videooverlaysoc_core_icmp_ip_port_source_payload_error;
assign soc_videooverlaysoc_core_icmp_rx_sink_sink_param_length = soc_videooverlaysoc_core_icmp_ip_port_source_param_length;
assign soc_videooverlaysoc_core_icmp_rx_sink_sink_param_protocol = soc_videooverlaysoc_core_icmp_ip_port_source_param_protocol;
assign soc_videooverlaysoc_core_icmp_rx_sink_sink_param_ip_address = soc_videooverlaysoc_core_icmp_ip_port_source_param_ip_address;
assign soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_valid = soc_videooverlaysoc_core_icmp_tx_sink_valid;
assign soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_last = soc_videooverlaysoc_core_icmp_tx_sink_last;
assign soc_videooverlaysoc_core_icmp_tx_sink_ready = soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_ready;
assign soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_msgtype = soc_videooverlaysoc_core_icmp_tx_sink_param_msgtype;
assign soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_code = soc_videooverlaysoc_core_icmp_tx_sink_param_code;
assign soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_checksum = soc_videooverlaysoc_core_icmp_tx_sink_param_checksum;
assign soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_quench = soc_videooverlaysoc_core_icmp_tx_sink_param_quench;
assign soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_payload_data = soc_videooverlaysoc_core_icmp_tx_sink_payload_data;
always @(*) begin
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header <= 64'd0;
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header[31:16] <= {soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_checksum[7:0], soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_checksum[15:8]};
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header[15:8] <= {soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_code[7:0]};
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header[7:0] <= {soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_msgtype[7:0]};
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header[63:32] <= {soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_quench[7:0], soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_quench[15:8], soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_quench[23:16], soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_param_quench[31:24]};
end
assign soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_payload_error = soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_payload_error;
always @(*) begin
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter_ce <= 1'd0;
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_valid <= 1'd0;
	vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_next_state <= 2'd0;
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_last <= 1'd0;
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_load <= 1'd0;
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_shift <= 1'd0;
	vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_next_state <= vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_state;
	case (vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_valid <= 1'd1;
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_last <= 1'd0;
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_payload_data <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header_reg[15:8];
			if ((soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_valid & soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_ready)) begin
				soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_shift <= 1'd1;
				soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter_ce <= 1'd1;
				if ((soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter == 3'd6)) begin
					vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_valid <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_valid;
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_last <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_last;
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_payload_data <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_payload_data;
			if ((soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_valid & soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_ready)) begin
				soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_ready <= 1'd1;
				if (soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_last) begin
					vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_valid) begin
				soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_sink_ready <= 1'd0;
				soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_valid <= 1'd1;
				soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_last <= 1'd0;
				soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_payload_data <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header[7:0];
				if ((soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_valid & soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_ready)) begin
					soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_load <= 1'd1;
					vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_next_state <= 1'd1;
				end
			end
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_core_icmp_tx_source_valid <= 1'd0;
	soc_videooverlaysoc_core_icmp_tx_source_first <= 1'd0;
	soc_videooverlaysoc_core_icmp_tx_source_last <= 1'd0;
	soc_videooverlaysoc_core_icmp_tx_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_ready <= 1'd0;
	soc_videooverlaysoc_core_icmp_tx_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_icmp_tx_source_param_length <= 16'd0;
	soc_videooverlaysoc_core_icmp_tx_source_param_protocol <= 8'd0;
	soc_videooverlaysoc_core_icmp_tx_source_param_ip_address <= 32'd0;
	vns_clockdomainsrenamer1_liteethicmptx_fsm_next_state <= 1'd0;
	vns_clockdomainsrenamer1_liteethicmptx_fsm_next_state <= vns_clockdomainsrenamer1_liteethicmptx_fsm_state;
	case (vns_clockdomainsrenamer1_liteethicmptx_fsm_state)
		1'd1: begin
			soc_videooverlaysoc_core_icmp_tx_source_valid <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_valid;
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_ready <= soc_videooverlaysoc_core_icmp_tx_source_ready;
			soc_videooverlaysoc_core_icmp_tx_source_first <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_first;
			soc_videooverlaysoc_core_icmp_tx_source_last <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_last;
			soc_videooverlaysoc_core_icmp_tx_source_payload_data <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_payload_data;
			soc_videooverlaysoc_core_icmp_tx_source_payload_error <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_payload_error;
			soc_videooverlaysoc_core_icmp_tx_source_param_length <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_param_length;
			soc_videooverlaysoc_core_icmp_tx_source_param_protocol <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_param_protocol;
			soc_videooverlaysoc_core_icmp_tx_source_param_ip_address <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_param_ip_address;
			soc_videooverlaysoc_core_icmp_tx_source_param_length <= (soc_videooverlaysoc_core_icmp_tx_sink_param_length + 4'd8);
			soc_videooverlaysoc_core_icmp_tx_source_param_protocol <= 1'd1;
			soc_videooverlaysoc_core_icmp_tx_source_param_ip_address <= soc_videooverlaysoc_core_icmp_tx_sink_param_ip_address;
			if (((soc_videooverlaysoc_core_icmp_tx_source_valid & soc_videooverlaysoc_core_icmp_tx_source_last) & soc_videooverlaysoc_core_icmp_tx_source_ready)) begin
				vns_clockdomainsrenamer1_liteethicmptx_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_ready <= 1'd1;
			if (soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_valid) begin
				soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_source_ready <= 1'd0;
				vns_clockdomainsrenamer1_liteethicmptx_fsm_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_valid = soc_videooverlaysoc_core_icmp_rx_sink_sink_valid;
assign soc_videooverlaysoc_core_icmp_rx_sink_sink_ready = soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_ready;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_first = soc_videooverlaysoc_core_icmp_rx_sink_sink_first;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_last = soc_videooverlaysoc_core_icmp_rx_sink_sink_last;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_payload_data = soc_videooverlaysoc_core_icmp_rx_sink_sink_payload_data;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_payload_error = soc_videooverlaysoc_core_icmp_rx_sink_sink_payload_error;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_param_length = soc_videooverlaysoc_core_icmp_rx_sink_sink_param_length;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_param_protocol = soc_videooverlaysoc_core_icmp_rx_sink_sink_param_protocol;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_param_ip_address = soc_videooverlaysoc_core_icmp_rx_sink_sink_param_ip_address;
assign soc_videooverlaysoc_core_icmp_rx_source_source_last = soc_videooverlaysoc_core_icmp_rx_depacketizer_source_last;
assign soc_videooverlaysoc_core_icmp_rx_source_source_param_msgtype = soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_msgtype;
assign soc_videooverlaysoc_core_icmp_rx_source_source_param_code = soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_code;
assign soc_videooverlaysoc_core_icmp_rx_source_source_param_checksum = soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_checksum;
assign soc_videooverlaysoc_core_icmp_rx_source_source_param_quench = soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_quench;
assign soc_videooverlaysoc_core_icmp_rx_source_source_param_ip_address = soc_videooverlaysoc_core_icmp_rx_sink_sink_param_ip_address;
assign soc_videooverlaysoc_core_icmp_rx_source_source_param_length = (soc_videooverlaysoc_core_icmp_rx_sink_sink_param_length - 4'd8);
assign soc_videooverlaysoc_core_icmp_rx_source_source_payload_data = soc_videooverlaysoc_core_icmp_rx_depacketizer_source_payload_data;
assign soc_videooverlaysoc_core_icmp_rx_source_source_payload_error = soc_videooverlaysoc_core_icmp_rx_depacketizer_source_payload_error;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_header = soc_videooverlaysoc_core_icmp_rx_depacketizer_header_reg;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_source_payload_error = soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_payload_error;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_source_last = (soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_last | soc_videooverlaysoc_core_icmp_rx_depacketizer_no_payload);
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_source_payload_data = soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_payload_data;
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_checksum = {vns_slice_proxy61[7:0], vns_slice_proxy60[15:8]};
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_code = {vns_slice_proxy62[7:0]};
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_msgtype = {vns_slice_proxy63[7:0]};
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_source_param_quench = {vns_slice_proxy67[7:0], vns_slice_proxy66[15:8], vns_slice_proxy65[23:16], vns_slice_proxy64[31:24]};
always @(*) begin
	soc_videooverlaysoc_core_icmp_rx_depacketizer_counter_ce <= 1'd0;
	soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_icmp_rx_depacketizer_source_valid <= 1'd0;
	soc_videooverlaysoc_core_icmp_rx_depacketizer_shift <= 1'd0;
	soc_videooverlaysoc_core_icmp_rx_depacketizer_counter_reset <= 1'd0;
	vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_next_state <= 2'd0;
	vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_next_state <= vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_state;
	case (vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_ready <= 1'd1;
			if (soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_valid) begin
				soc_videooverlaysoc_core_icmp_rx_depacketizer_counter_ce <= 1'd1;
				soc_videooverlaysoc_core_icmp_rx_depacketizer_shift <= 1'd1;
				if ((soc_videooverlaysoc_core_icmp_rx_depacketizer_counter == 3'd6)) begin
					vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_ready <= soc_videooverlaysoc_core_icmp_rx_depacketizer_source_ready;
			soc_videooverlaysoc_core_icmp_rx_depacketizer_source_valid <= (soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_valid | soc_videooverlaysoc_core_icmp_rx_depacketizer_no_payload);
			if (((soc_videooverlaysoc_core_icmp_rx_depacketizer_source_valid & soc_videooverlaysoc_core_icmp_rx_depacketizer_source_ready) & soc_videooverlaysoc_core_icmp_rx_depacketizer_source_last)) begin
				vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_icmp_rx_depacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_valid) begin
				soc_videooverlaysoc_core_icmp_rx_depacketizer_shift <= 1'd1;
				vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_icmp_rx_depacketizer_is_el = ((~(vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_state == 2'd2)) & (vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_next_state == 2'd2));
always @(*) begin
	soc_videooverlaysoc_core_icmp_rx_source_source_valid <= 1'd0;
	soc_videooverlaysoc_core_icmp_rx_depacketizer_source_ready <= 1'd0;
	vns_clockdomainsrenamer1_liteethicmprx_fsm_next_state <= 2'd0;
	vns_clockdomainsrenamer1_liteethicmprx_fsm_next_state <= vns_clockdomainsrenamer1_liteethicmprx_fsm_state;
	case (vns_clockdomainsrenamer1_liteethicmprx_fsm_state)
		1'd1: begin
			if (soc_videooverlaysoc_core_icmp_rx_valid) begin
				vns_clockdomainsrenamer1_liteethicmprx_fsm_next_state <= 2'd2;
			end else begin
				vns_clockdomainsrenamer1_liteethicmprx_fsm_next_state <= 2'd3;
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_icmp_rx_source_source_valid <= soc_videooverlaysoc_core_icmp_rx_depacketizer_source_valid;
			soc_videooverlaysoc_core_icmp_rx_depacketizer_source_ready <= soc_videooverlaysoc_core_icmp_rx_source_source_ready;
			if (((soc_videooverlaysoc_core_icmp_rx_source_source_valid & soc_videooverlaysoc_core_icmp_rx_source_source_last) & soc_videooverlaysoc_core_icmp_rx_source_source_ready)) begin
				vns_clockdomainsrenamer1_liteethicmprx_fsm_next_state <= 1'd0;
			end
		end
		2'd3: begin
			soc_videooverlaysoc_core_icmp_rx_depacketizer_source_ready <= 1'd1;
			if (((soc_videooverlaysoc_core_icmp_rx_depacketizer_source_valid & soc_videooverlaysoc_core_icmp_rx_depacketizer_source_last) & soc_videooverlaysoc_core_icmp_rx_depacketizer_source_ready)) begin
				vns_clockdomainsrenamer1_liteethicmprx_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_icmp_rx_depacketizer_source_ready <= 1'd1;
			if (soc_videooverlaysoc_core_icmp_rx_depacketizer_source_valid) begin
				soc_videooverlaysoc_core_icmp_rx_depacketizer_source_ready <= 1'd0;
				vns_clockdomainsrenamer1_liteethicmprx_fsm_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_valid = soc_videooverlaysoc_core_icmp_echo_sink_sink_valid;
assign soc_videooverlaysoc_core_icmp_echo_sink_sink_ready = soc_videooverlaysoc_core_icmp_echo_buffer_sink_ready;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_first = soc_videooverlaysoc_core_icmp_echo_sink_sink_first;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_last = soc_videooverlaysoc_core_icmp_echo_sink_sink_last;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_payload_data = soc_videooverlaysoc_core_icmp_echo_sink_sink_payload_data;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_payload_error = soc_videooverlaysoc_core_icmp_echo_sink_sink_payload_error;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_checksum = soc_videooverlaysoc_core_icmp_echo_sink_sink_param_checksum;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_code = soc_videooverlaysoc_core_icmp_echo_sink_sink_param_code;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_msgtype = soc_videooverlaysoc_core_icmp_echo_sink_sink_param_msgtype;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_quench = soc_videooverlaysoc_core_icmp_echo_sink_sink_param_quench;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_ip_address = soc_videooverlaysoc_core_icmp_echo_sink_sink_param_ip_address;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_length = soc_videooverlaysoc_core_icmp_echo_sink_sink_param_length;
assign soc_videooverlaysoc_core_icmp_echo_source_source_valid = soc_videooverlaysoc_core_icmp_echo_buffer_source_valid;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_ready = soc_videooverlaysoc_core_icmp_echo_source_source_ready;
assign soc_videooverlaysoc_core_icmp_echo_source_source_first = soc_videooverlaysoc_core_icmp_echo_buffer_source_first;
assign soc_videooverlaysoc_core_icmp_echo_source_source_last = soc_videooverlaysoc_core_icmp_echo_buffer_source_last;
assign soc_videooverlaysoc_core_icmp_echo_source_source_payload_data = soc_videooverlaysoc_core_icmp_echo_buffer_source_payload_data;
assign soc_videooverlaysoc_core_icmp_echo_source_source_payload_error = soc_videooverlaysoc_core_icmp_echo_buffer_source_payload_error;
assign soc_videooverlaysoc_core_icmp_echo_source_source_param_code = soc_videooverlaysoc_core_icmp_echo_buffer_source_param_code;
assign soc_videooverlaysoc_core_icmp_echo_source_source_param_quench = soc_videooverlaysoc_core_icmp_echo_buffer_source_param_quench;
assign soc_videooverlaysoc_core_icmp_echo_source_source_param_ip_address = soc_videooverlaysoc_core_icmp_echo_buffer_source_param_ip_address;
assign soc_videooverlaysoc_core_icmp_echo_source_source_param_length = soc_videooverlaysoc_core_icmp_echo_buffer_source_param_length;
always @(*) begin
	soc_videooverlaysoc_core_icmp_echo_source_source_param_msgtype <= 8'd0;
	soc_videooverlaysoc_core_icmp_echo_source_source_param_msgtype <= soc_videooverlaysoc_core_icmp_echo_buffer_source_param_msgtype;
	soc_videooverlaysoc_core_icmp_echo_source_source_param_msgtype <= 1'd0;
end
always @(*) begin
	soc_videooverlaysoc_core_icmp_echo_source_source_param_checksum <= 16'd0;
	soc_videooverlaysoc_core_icmp_echo_source_source_param_checksum <= soc_videooverlaysoc_core_icmp_echo_buffer_source_param_checksum;
	soc_videooverlaysoc_core_icmp_echo_source_source_param_checksum <= (~((~soc_videooverlaysoc_core_icmp_echo_buffer_source_param_checksum) - 12'd2048));
end
assign soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_din = {soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_last, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_first, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_length, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_ip_address, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_quench, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_msgtype, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_code, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_checksum, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_payload_error, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_payload_data};
assign {soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_last, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_first, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_length, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_ip_address, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_quench, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_msgtype, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_code, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_checksum, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_payload_error, soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_payload_data} = soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_dout;
assign soc_videooverlaysoc_core_icmp_echo_buffer_sink_ready = soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_writable;
assign soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_we = soc_videooverlaysoc_core_icmp_echo_buffer_sink_valid;
assign soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_first = soc_videooverlaysoc_core_icmp_echo_buffer_sink_first;
assign soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_last = soc_videooverlaysoc_core_icmp_echo_buffer_sink_last;
assign soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_payload_data = soc_videooverlaysoc_core_icmp_echo_buffer_sink_payload_data;
assign soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_payload_error = soc_videooverlaysoc_core_icmp_echo_buffer_sink_payload_error;
assign soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_checksum = soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_checksum;
assign soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_code = soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_code;
assign soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_msgtype = soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_msgtype;
assign soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_quench = soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_quench;
assign soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_ip_address = soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_ip_address;
assign soc_videooverlaysoc_core_icmp_echo_buffer_fifo_in_param_length = soc_videooverlaysoc_core_icmp_echo_buffer_sink_param_length;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_valid = soc_videooverlaysoc_core_icmp_echo_buffer_readable;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_first = soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_first;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_last = soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_last;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_payload_data = soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_payload_data;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_payload_error = soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_payload_error;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_param_checksum = soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_checksum;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_param_code = soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_code;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_param_msgtype = soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_msgtype;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_param_quench = soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_quench;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_param_ip_address = soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_ip_address;
assign soc_videooverlaysoc_core_icmp_echo_buffer_source_param_length = soc_videooverlaysoc_core_icmp_echo_buffer_fifo_out_param_length;
assign soc_videooverlaysoc_core_icmp_echo_buffer_re = soc_videooverlaysoc_core_icmp_echo_buffer_source_ready;
assign soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_re = (soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_readable & ((~soc_videooverlaysoc_core_icmp_echo_buffer_readable) | soc_videooverlaysoc_core_icmp_echo_buffer_re));
assign soc_videooverlaysoc_core_icmp_echo_buffer_level1 = (soc_videooverlaysoc_core_icmp_echo_buffer_level0 + soc_videooverlaysoc_core_icmp_echo_buffer_readable);
always @(*) begin
	soc_videooverlaysoc_core_icmp_echo_buffer_wrport_adr <= 7'd0;
	if (soc_videooverlaysoc_core_icmp_echo_buffer_replace) begin
		soc_videooverlaysoc_core_icmp_echo_buffer_wrport_adr <= (soc_videooverlaysoc_core_icmp_echo_buffer_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_core_icmp_echo_buffer_wrport_adr <= soc_videooverlaysoc_core_icmp_echo_buffer_produce;
	end
end
assign soc_videooverlaysoc_core_icmp_echo_buffer_wrport_dat_w = soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_din;
assign soc_videooverlaysoc_core_icmp_echo_buffer_wrport_we = (soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_we & (soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_writable | soc_videooverlaysoc_core_icmp_echo_buffer_replace));
assign soc_videooverlaysoc_core_icmp_echo_buffer_do_read = (soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_readable & soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_re);
assign soc_videooverlaysoc_core_icmp_echo_buffer_rdport_adr = soc_videooverlaysoc_core_icmp_echo_buffer_consume;
assign soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_dout = soc_videooverlaysoc_core_icmp_echo_buffer_rdport_dat_r;
assign soc_videooverlaysoc_core_icmp_echo_buffer_rdport_re = soc_videooverlaysoc_core_icmp_echo_buffer_do_read;
assign soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_writable = (soc_videooverlaysoc_core_icmp_echo_buffer_level0 != 8'd128);
assign soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_readable = (soc_videooverlaysoc_core_icmp_echo_buffer_level0 != 1'd0);
assign soc_videooverlaysoc_core_ip_port_sink_valid = soc_videooverlaysoc_core_tx_source_valid;
assign soc_videooverlaysoc_core_tx_source_ready = soc_videooverlaysoc_core_ip_port_sink_ready;
assign soc_videooverlaysoc_core_ip_port_sink_first = soc_videooverlaysoc_core_tx_source_first;
assign soc_videooverlaysoc_core_ip_port_sink_last = soc_videooverlaysoc_core_tx_source_last;
assign soc_videooverlaysoc_core_ip_port_sink_payload_data = soc_videooverlaysoc_core_tx_source_payload_data;
assign soc_videooverlaysoc_core_ip_port_sink_payload_error = soc_videooverlaysoc_core_tx_source_payload_error;
assign soc_videooverlaysoc_core_ip_port_sink_param_length = soc_videooverlaysoc_core_tx_source_param_length;
assign soc_videooverlaysoc_core_ip_port_sink_param_protocol = soc_videooverlaysoc_core_tx_source_param_protocol;
assign soc_videooverlaysoc_core_ip_port_sink_param_ip_address = soc_videooverlaysoc_core_tx_source_param_ip_address;
assign soc_videooverlaysoc_core_sink_sink_valid = soc_videooverlaysoc_core_ip_port_source_valid;
assign soc_videooverlaysoc_core_ip_port_source_ready = soc_videooverlaysoc_core_sink_sink_ready;
assign soc_videooverlaysoc_core_sink_sink_first = soc_videooverlaysoc_core_ip_port_source_first;
assign soc_videooverlaysoc_core_sink_sink_last = soc_videooverlaysoc_core_ip_port_source_last;
assign soc_videooverlaysoc_core_sink_sink_payload_data = soc_videooverlaysoc_core_ip_port_source_payload_data;
assign soc_videooverlaysoc_core_sink_sink_payload_error = soc_videooverlaysoc_core_ip_port_source_payload_error;
assign soc_videooverlaysoc_core_sink_sink_param_length = soc_videooverlaysoc_core_ip_port_source_param_length;
assign soc_videooverlaysoc_core_sink_sink_param_protocol = soc_videooverlaysoc_core_ip_port_source_param_protocol;
assign soc_videooverlaysoc_core_sink_sink_param_ip_address = soc_videooverlaysoc_core_ip_port_source_param_ip_address;
assign soc_videooverlaysoc_core_tx_sink_valid = soc_videooverlaysoc_core_crossbar_source_valid;
assign soc_videooverlaysoc_core_crossbar_source_ready = soc_videooverlaysoc_core_tx_sink_ready;
assign soc_videooverlaysoc_core_tx_sink_first = soc_videooverlaysoc_core_crossbar_source_first;
assign soc_videooverlaysoc_core_tx_sink_last = soc_videooverlaysoc_core_crossbar_source_last;
assign soc_videooverlaysoc_core_tx_sink_payload_data = soc_videooverlaysoc_core_crossbar_source_payload_data;
assign soc_videooverlaysoc_core_tx_sink_payload_error = soc_videooverlaysoc_core_crossbar_source_payload_error;
assign soc_videooverlaysoc_core_tx_sink_param_src_port = soc_videooverlaysoc_core_crossbar_source_param_src_port;
assign soc_videooverlaysoc_core_tx_sink_param_dst_port = soc_videooverlaysoc_core_crossbar_source_param_dst_port;
assign soc_videooverlaysoc_core_tx_sink_param_ip_address = soc_videooverlaysoc_core_crossbar_source_param_ip_address;
assign soc_videooverlaysoc_core_tx_sink_param_length = soc_videooverlaysoc_core_crossbar_source_param_length;
assign soc_videooverlaysoc_core_crossbar_sink_valid = soc_videooverlaysoc_core_source_source_valid;
assign soc_videooverlaysoc_core_source_source_ready = soc_videooverlaysoc_core_crossbar_sink_ready;
assign soc_videooverlaysoc_core_crossbar_sink_first = soc_videooverlaysoc_core_source_source_first;
assign soc_videooverlaysoc_core_crossbar_sink_last = soc_videooverlaysoc_core_source_source_last;
assign soc_videooverlaysoc_core_crossbar_sink_payload_data = soc_videooverlaysoc_core_source_source_payload_data;
assign soc_videooverlaysoc_core_crossbar_sink_payload_error = soc_videooverlaysoc_core_source_source_payload_error;
assign soc_videooverlaysoc_core_crossbar_sink_param_src_port = soc_videooverlaysoc_core_source_source_param_src_port;
assign soc_videooverlaysoc_core_crossbar_sink_param_dst_port = soc_videooverlaysoc_core_source_source_param_dst_port;
assign soc_videooverlaysoc_core_crossbar_sink_param_ip_address = soc_videooverlaysoc_core_source_source_param_ip_address;
assign soc_videooverlaysoc_core_crossbar_sink_param_length = soc_videooverlaysoc_core_source_source_param_length;
assign soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_valid = soc_videooverlaysoc_core_tx_sink_valid;
assign soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_last = soc_videooverlaysoc_core_tx_sink_last;
assign soc_videooverlaysoc_core_tx_sink_ready = soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_ready;
assign soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_src_port = soc_videooverlaysoc_core_tx_sink_param_src_port;
assign soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_dst_port = soc_videooverlaysoc_core_tx_sink_param_dst_port;
assign soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_length = (soc_videooverlaysoc_core_tx_sink_param_length + 4'd8);
assign soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_checksum = 1'd0;
assign soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_payload_data = soc_videooverlaysoc_core_tx_sink_payload_data;
always @(*) begin
	soc_videooverlaysoc_core_tx_liteethudppacketizer_header <= 64'd0;
	soc_videooverlaysoc_core_tx_liteethudppacketizer_header[63:48] <= {soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_checksum[7:0], soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_checksum[15:8]};
	soc_videooverlaysoc_core_tx_liteethudppacketizer_header[31:16] <= {soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_dst_port[7:0], soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_dst_port[15:8]};
	soc_videooverlaysoc_core_tx_liteethudppacketizer_header[47:32] <= {soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_length[7:0], soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_length[15:8]};
	soc_videooverlaysoc_core_tx_liteethudppacketizer_header[15:0] <= {soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_src_port[7:0], soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_src_port[15:8]};
end
assign soc_videooverlaysoc_core_tx_liteethudppacketizer_source_payload_error = soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_payload_error;
always @(*) begin
	soc_videooverlaysoc_core_tx_liteethudppacketizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_tx_liteethudppacketizer_counter_ce <= 1'd0;
	soc_videooverlaysoc_core_tx_liteethudppacketizer_source_valid <= 1'd0;
	vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_next_state <= 2'd0;
	soc_videooverlaysoc_core_tx_liteethudppacketizer_source_last <= 1'd0;
	soc_videooverlaysoc_core_tx_liteethudppacketizer_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_tx_liteethudppacketizer_load <= 1'd0;
	soc_videooverlaysoc_core_tx_liteethudppacketizer_shift <= 1'd0;
	vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_next_state <= vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_state;
	case (vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_core_tx_liteethudppacketizer_source_valid <= 1'd1;
			soc_videooverlaysoc_core_tx_liteethudppacketizer_source_last <= 1'd0;
			soc_videooverlaysoc_core_tx_liteethudppacketizer_source_payload_data <= soc_videooverlaysoc_core_tx_liteethudppacketizer_header_reg[15:8];
			if ((soc_videooverlaysoc_core_tx_liteethudppacketizer_source_valid & soc_videooverlaysoc_core_tx_liteethudppacketizer_source_ready)) begin
				soc_videooverlaysoc_core_tx_liteethudppacketizer_shift <= 1'd1;
				soc_videooverlaysoc_core_tx_liteethudppacketizer_counter_ce <= 1'd1;
				if ((soc_videooverlaysoc_core_tx_liteethudppacketizer_counter == 3'd6)) begin
					vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_tx_liteethudppacketizer_source_valid <= soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_valid;
			soc_videooverlaysoc_core_tx_liteethudppacketizer_source_last <= soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_last;
			soc_videooverlaysoc_core_tx_liteethudppacketizer_source_payload_data <= soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_payload_data;
			if ((soc_videooverlaysoc_core_tx_liteethudppacketizer_source_valid & soc_videooverlaysoc_core_tx_liteethudppacketizer_source_ready)) begin
				soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_ready <= 1'd1;
				if (soc_videooverlaysoc_core_tx_liteethudppacketizer_source_last) begin
					vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_tx_liteethudppacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_valid) begin
				soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_ready <= 1'd0;
				soc_videooverlaysoc_core_tx_liteethudppacketizer_source_valid <= 1'd1;
				soc_videooverlaysoc_core_tx_liteethudppacketizer_source_last <= 1'd0;
				soc_videooverlaysoc_core_tx_liteethudppacketizer_source_payload_data <= soc_videooverlaysoc_core_tx_liteethudppacketizer_header[7:0];
				if ((soc_videooverlaysoc_core_tx_liteethudppacketizer_source_valid & soc_videooverlaysoc_core_tx_liteethudppacketizer_source_ready)) begin
					soc_videooverlaysoc_core_tx_liteethudppacketizer_load <= 1'd1;
					vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_next_state <= 1'd1;
				end
			end
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_core_tx_source_valid <= 1'd0;
	soc_videooverlaysoc_core_tx_source_first <= 1'd0;
	soc_videooverlaysoc_core_tx_source_last <= 1'd0;
	soc_videooverlaysoc_core_tx_source_payload_data <= 8'd0;
	soc_videooverlaysoc_core_tx_liteethudppacketizer_source_ready <= 1'd0;
	soc_videooverlaysoc_core_tx_source_payload_error <= 1'd0;
	soc_videooverlaysoc_core_tx_source_param_length <= 16'd0;
	soc_videooverlaysoc_core_tx_source_param_protocol <= 8'd0;
	soc_videooverlaysoc_core_tx_source_param_ip_address <= 32'd0;
	vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_next_state <= 1'd0;
	vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_next_state <= vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_state;
	case (vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_state)
		1'd1: begin
			soc_videooverlaysoc_core_tx_source_valid <= soc_videooverlaysoc_core_tx_liteethudppacketizer_source_valid;
			soc_videooverlaysoc_core_tx_liteethudppacketizer_source_ready <= soc_videooverlaysoc_core_tx_source_ready;
			soc_videooverlaysoc_core_tx_source_first <= soc_videooverlaysoc_core_tx_liteethudppacketizer_source_first;
			soc_videooverlaysoc_core_tx_source_last <= soc_videooverlaysoc_core_tx_liteethudppacketizer_source_last;
			soc_videooverlaysoc_core_tx_source_payload_data <= soc_videooverlaysoc_core_tx_liteethudppacketizer_source_payload_data;
			soc_videooverlaysoc_core_tx_source_payload_error <= soc_videooverlaysoc_core_tx_liteethudppacketizer_source_payload_error;
			soc_videooverlaysoc_core_tx_source_param_length <= soc_videooverlaysoc_core_tx_liteethudppacketizer_source_param_length;
			soc_videooverlaysoc_core_tx_source_param_protocol <= soc_videooverlaysoc_core_tx_liteethudppacketizer_source_param_protocol;
			soc_videooverlaysoc_core_tx_source_param_ip_address <= soc_videooverlaysoc_core_tx_liteethudppacketizer_source_param_ip_address;
			soc_videooverlaysoc_core_tx_source_param_length <= soc_videooverlaysoc_core_tx_liteethudppacketizer_sink_param_length;
			soc_videooverlaysoc_core_tx_source_param_protocol <= 5'd17;
			soc_videooverlaysoc_core_tx_source_param_ip_address <= soc_videooverlaysoc_core_tx_sink_param_ip_address;
			if (((soc_videooverlaysoc_core_tx_source_valid & soc_videooverlaysoc_core_tx_source_last) & soc_videooverlaysoc_core_tx_source_ready)) begin
				vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_tx_liteethudppacketizer_source_ready <= 1'd1;
			if (soc_videooverlaysoc_core_tx_liteethudppacketizer_source_valid) begin
				soc_videooverlaysoc_core_tx_liteethudppacketizer_source_ready <= 1'd0;
				vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_depacketizer_sink_valid = soc_videooverlaysoc_core_sink_sink_valid;
assign soc_videooverlaysoc_core_sink_sink_ready = soc_videooverlaysoc_core_depacketizer_sink_ready;
assign soc_videooverlaysoc_core_depacketizer_sink_first = soc_videooverlaysoc_core_sink_sink_first;
assign soc_videooverlaysoc_core_depacketizer_sink_last = soc_videooverlaysoc_core_sink_sink_last;
assign soc_videooverlaysoc_core_depacketizer_sink_payload_data = soc_videooverlaysoc_core_sink_sink_payload_data;
assign soc_videooverlaysoc_core_depacketizer_sink_payload_error = soc_videooverlaysoc_core_sink_sink_payload_error;
assign soc_videooverlaysoc_core_depacketizer_sink_param_length = soc_videooverlaysoc_core_sink_sink_param_length;
assign soc_videooverlaysoc_core_depacketizer_sink_param_protocol = soc_videooverlaysoc_core_sink_sink_param_protocol;
assign soc_videooverlaysoc_core_depacketizer_sink_param_ip_address = soc_videooverlaysoc_core_sink_sink_param_ip_address;
assign soc_videooverlaysoc_core_source_source_last = soc_videooverlaysoc_core_depacketizer_source_last;
assign soc_videooverlaysoc_core_source_source_param_src_port = soc_videooverlaysoc_core_depacketizer_source_param_src_port;
assign soc_videooverlaysoc_core_source_source_param_dst_port = soc_videooverlaysoc_core_depacketizer_source_param_dst_port;
assign soc_videooverlaysoc_core_source_source_param_ip_address = soc_videooverlaysoc_core_sink_sink_param_ip_address;
assign soc_videooverlaysoc_core_source_source_param_length = (soc_videooverlaysoc_core_depacketizer_source_param_length - 4'd8);
assign soc_videooverlaysoc_core_source_source_payload_data = soc_videooverlaysoc_core_depacketizer_source_payload_data;
assign soc_videooverlaysoc_core_source_source_payload_error = soc_videooverlaysoc_core_depacketizer_source_payload_error;
assign soc_videooverlaysoc_core_depacketizer_header = soc_videooverlaysoc_core_depacketizer_header_reg;
assign soc_videooverlaysoc_core_depacketizer_source_payload_error = soc_videooverlaysoc_core_depacketizer_sink_payload_error;
assign soc_videooverlaysoc_core_depacketizer_source_last = (soc_videooverlaysoc_core_depacketizer_sink_last | soc_videooverlaysoc_core_depacketizer_no_payload);
assign soc_videooverlaysoc_core_depacketizer_source_payload_data = soc_videooverlaysoc_core_depacketizer_sink_payload_data;
assign soc_videooverlaysoc_core_depacketizer_source_param_checksum = {vns_slice_proxy69[7:0], vns_slice_proxy68[15:8]};
assign soc_videooverlaysoc_core_depacketizer_source_param_dst_port = {vns_slice_proxy71[7:0], vns_slice_proxy70[15:8]};
assign soc_videooverlaysoc_core_depacketizer_source_param_length = {vns_slice_proxy73[7:0], vns_slice_proxy72[15:8]};
assign soc_videooverlaysoc_core_depacketizer_source_param_src_port = {vns_slice_proxy75[7:0], vns_slice_proxy74[15:8]};
always @(*) begin
	soc_videooverlaysoc_core_depacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_core_depacketizer_source_valid <= 1'd0;
	soc_videooverlaysoc_core_depacketizer_shift <= 1'd0;
	vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_next_state <= 2'd0;
	soc_videooverlaysoc_core_depacketizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_core_depacketizer_counter_ce <= 1'd0;
	vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_next_state <= vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_state;
	case (vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_core_depacketizer_sink_ready <= 1'd1;
			if (soc_videooverlaysoc_core_depacketizer_sink_valid) begin
				soc_videooverlaysoc_core_depacketizer_counter_ce <= 1'd1;
				soc_videooverlaysoc_core_depacketizer_shift <= 1'd1;
				if ((soc_videooverlaysoc_core_depacketizer_counter == 3'd6)) begin
					vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_depacketizer_sink_ready <= soc_videooverlaysoc_core_depacketizer_source_ready;
			soc_videooverlaysoc_core_depacketizer_source_valid <= (soc_videooverlaysoc_core_depacketizer_sink_valid | soc_videooverlaysoc_core_depacketizer_no_payload);
			if (((soc_videooverlaysoc_core_depacketizer_source_valid & soc_videooverlaysoc_core_depacketizer_source_ready) & soc_videooverlaysoc_core_depacketizer_source_last)) begin
				vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_depacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_core_depacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_core_depacketizer_sink_valid) begin
				soc_videooverlaysoc_core_depacketizer_shift <= 1'd1;
				vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_core_depacketizer_is_el = ((~(vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_state == 2'd2)) & (vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_next_state == 2'd2));
always @(*) begin
	vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_next_state <= 2'd0;
	soc_videooverlaysoc_core_source_source_valid <= 1'd0;
	soc_videooverlaysoc_core_depacketizer_source_ready <= 1'd0;
	vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_next_state <= vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_state;
	case (vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_state)
		1'd1: begin
			if (soc_videooverlaysoc_core_valid) begin
				vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_next_state <= 2'd2;
			end else begin
				vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_next_state <= 2'd3;
			end
		end
		2'd2: begin
			soc_videooverlaysoc_core_source_source_valid <= soc_videooverlaysoc_core_depacketizer_source_valid;
			soc_videooverlaysoc_core_depacketizer_source_ready <= soc_videooverlaysoc_core_source_source_ready;
			if (((soc_videooverlaysoc_core_source_source_valid & soc_videooverlaysoc_core_source_source_last) & soc_videooverlaysoc_core_source_source_ready)) begin
				vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_next_state <= 1'd0;
			end
		end
		2'd3: begin
			soc_videooverlaysoc_core_depacketizer_source_ready <= 1'd1;
			if (((soc_videooverlaysoc_core_depacketizer_source_valid & soc_videooverlaysoc_core_depacketizer_source_last) & soc_videooverlaysoc_core_depacketizer_source_ready)) begin
				vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_core_depacketizer_source_ready <= 1'd1;
			if (soc_videooverlaysoc_core_depacketizer_source_valid) begin
				soc_videooverlaysoc_core_depacketizer_source_ready <= 1'd0;
				vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_packet_tx_cdc_sink_valid = soc_videooverlaysoc_packet_user_port_sink_valid;
assign soc_videooverlaysoc_packet_user_port_sink_ready = soc_videooverlaysoc_packet_tx_cdc_sink_ready;
assign soc_videooverlaysoc_packet_tx_cdc_sink_first = soc_videooverlaysoc_packet_user_port_sink_first;
assign soc_videooverlaysoc_packet_tx_cdc_sink_last = soc_videooverlaysoc_packet_user_port_sink_last;
assign soc_videooverlaysoc_packet_tx_cdc_sink_payload_data = soc_videooverlaysoc_packet_user_port_sink_payload_data;
assign soc_videooverlaysoc_packet_tx_cdc_sink_payload_error = soc_videooverlaysoc_packet_user_port_sink_payload_error;
assign soc_videooverlaysoc_packet_tx_cdc_sink_param_src_port = soc_videooverlaysoc_packet_user_port_sink_param_src_port;
assign soc_videooverlaysoc_packet_tx_cdc_sink_param_dst_port = soc_videooverlaysoc_packet_user_port_sink_param_dst_port;
assign soc_videooverlaysoc_packet_tx_cdc_sink_param_ip_address = soc_videooverlaysoc_packet_user_port_sink_param_ip_address;
assign soc_videooverlaysoc_packet_tx_cdc_sink_param_length = soc_videooverlaysoc_packet_user_port_sink_param_length;
assign soc_videooverlaysoc_packet_tx_converter_sink_valid = soc_videooverlaysoc_packet_tx_cdc_source_valid;
assign soc_videooverlaysoc_packet_tx_cdc_source_ready = soc_videooverlaysoc_packet_tx_converter_sink_ready;
assign soc_videooverlaysoc_packet_tx_converter_sink_first = soc_videooverlaysoc_packet_tx_cdc_source_first;
assign soc_videooverlaysoc_packet_tx_converter_sink_last = soc_videooverlaysoc_packet_tx_cdc_source_last;
assign soc_videooverlaysoc_packet_tx_converter_sink_payload_data = soc_videooverlaysoc_packet_tx_cdc_source_payload_data;
assign soc_videooverlaysoc_packet_tx_converter_sink_payload_error = soc_videooverlaysoc_packet_tx_cdc_source_payload_error;
assign soc_videooverlaysoc_packet_tx_converter_sink_param_src_port = soc_videooverlaysoc_packet_tx_cdc_source_param_src_port;
assign soc_videooverlaysoc_packet_tx_converter_sink_param_dst_port = soc_videooverlaysoc_packet_tx_cdc_source_param_dst_port;
assign soc_videooverlaysoc_packet_tx_converter_sink_param_ip_address = soc_videooverlaysoc_packet_tx_cdc_source_param_ip_address;
assign soc_videooverlaysoc_packet_tx_converter_sink_param_length = soc_videooverlaysoc_packet_tx_cdc_source_param_length;
assign soc_videooverlaysoc_packet_internal_port_sink_valid = soc_videooverlaysoc_packet_tx_converter_source_valid;
assign soc_videooverlaysoc_packet_tx_converter_source_ready = soc_videooverlaysoc_packet_internal_port_sink_ready;
assign soc_videooverlaysoc_packet_internal_port_sink_first = soc_videooverlaysoc_packet_tx_converter_source_first;
assign soc_videooverlaysoc_packet_internal_port_sink_last = soc_videooverlaysoc_packet_tx_converter_source_last;
assign soc_videooverlaysoc_packet_internal_port_sink_payload_data = soc_videooverlaysoc_packet_tx_converter_source_payload_data;
assign soc_videooverlaysoc_packet_internal_port_sink_payload_error = soc_videooverlaysoc_packet_tx_converter_source_payload_error;
assign soc_videooverlaysoc_packet_internal_port_sink_param_src_port = soc_videooverlaysoc_packet_tx_converter_source_param_src_port;
assign soc_videooverlaysoc_packet_internal_port_sink_param_dst_port = soc_videooverlaysoc_packet_tx_converter_source_param_dst_port;
assign soc_videooverlaysoc_packet_internal_port_sink_param_ip_address = soc_videooverlaysoc_packet_tx_converter_source_param_ip_address;
assign soc_videooverlaysoc_packet_internal_port_sink_param_length = soc_videooverlaysoc_packet_tx_converter_source_param_length;
assign soc_videooverlaysoc_packet_rx_converter_sink_valid = soc_videooverlaysoc_packet_internal_port_source_valid;
assign soc_videooverlaysoc_packet_internal_port_source_ready = soc_videooverlaysoc_packet_rx_converter_sink_ready;
assign soc_videooverlaysoc_packet_rx_converter_sink_first = soc_videooverlaysoc_packet_internal_port_source_first;
assign soc_videooverlaysoc_packet_rx_converter_sink_last = soc_videooverlaysoc_packet_internal_port_source_last;
assign soc_videooverlaysoc_packet_rx_converter_sink_payload_data = soc_videooverlaysoc_packet_internal_port_source_payload_data;
assign soc_videooverlaysoc_packet_rx_converter_sink_payload_error = soc_videooverlaysoc_packet_internal_port_source_payload_error;
assign soc_videooverlaysoc_packet_rx_converter_sink_param_src_port = soc_videooverlaysoc_packet_internal_port_source_param_src_port;
assign soc_videooverlaysoc_packet_rx_converter_sink_param_dst_port = soc_videooverlaysoc_packet_internal_port_source_param_dst_port;
assign soc_videooverlaysoc_packet_rx_converter_sink_param_ip_address = soc_videooverlaysoc_packet_internal_port_source_param_ip_address;
assign soc_videooverlaysoc_packet_rx_converter_sink_param_length = soc_videooverlaysoc_packet_internal_port_source_param_length;
assign soc_videooverlaysoc_packet_rx_cdc_sink_valid = soc_videooverlaysoc_packet_rx_converter_source_valid;
assign soc_videooverlaysoc_packet_rx_converter_source_ready = soc_videooverlaysoc_packet_rx_cdc_sink_ready;
assign soc_videooverlaysoc_packet_rx_cdc_sink_first = soc_videooverlaysoc_packet_rx_converter_source_first;
assign soc_videooverlaysoc_packet_rx_cdc_sink_last = soc_videooverlaysoc_packet_rx_converter_source_last;
assign soc_videooverlaysoc_packet_rx_cdc_sink_payload_data = soc_videooverlaysoc_packet_rx_converter_source_payload_data;
assign soc_videooverlaysoc_packet_rx_cdc_sink_payload_error = soc_videooverlaysoc_packet_rx_converter_source_payload_error;
assign soc_videooverlaysoc_packet_rx_cdc_sink_param_src_port = soc_videooverlaysoc_packet_rx_converter_source_param_src_port;
assign soc_videooverlaysoc_packet_rx_cdc_sink_param_dst_port = soc_videooverlaysoc_packet_rx_converter_source_param_dst_port;
assign soc_videooverlaysoc_packet_rx_cdc_sink_param_ip_address = soc_videooverlaysoc_packet_rx_converter_source_param_ip_address;
assign soc_videooverlaysoc_packet_rx_cdc_sink_param_length = soc_videooverlaysoc_packet_rx_converter_source_param_length;
assign soc_videooverlaysoc_packet_user_port_source_valid = soc_videooverlaysoc_packet_rx_cdc_source_valid;
assign soc_videooverlaysoc_packet_rx_cdc_source_ready = soc_videooverlaysoc_packet_user_port_source_ready;
assign soc_videooverlaysoc_packet_user_port_source_first = soc_videooverlaysoc_packet_rx_cdc_source_first;
assign soc_videooverlaysoc_packet_user_port_source_last = soc_videooverlaysoc_packet_rx_cdc_source_last;
assign soc_videooverlaysoc_packet_user_port_source_payload_data = soc_videooverlaysoc_packet_rx_cdc_source_payload_data;
assign soc_videooverlaysoc_packet_user_port_source_payload_error = soc_videooverlaysoc_packet_rx_cdc_source_payload_error;
assign soc_videooverlaysoc_packet_user_port_source_param_src_port = soc_videooverlaysoc_packet_rx_cdc_source_param_src_port;
assign soc_videooverlaysoc_packet_user_port_source_param_dst_port = soc_videooverlaysoc_packet_rx_cdc_source_param_dst_port;
assign soc_videooverlaysoc_packet_user_port_source_param_ip_address = soc_videooverlaysoc_packet_rx_cdc_source_param_ip_address;
assign soc_videooverlaysoc_packet_user_port_source_param_length = soc_videooverlaysoc_packet_rx_cdc_source_param_length;
always @(*) begin
	vns_clockdomainsrenamer1_liteethudp_sel <= 1'd0;
	case (soc_videooverlaysoc_core_crossbar_sink_param_dst_port)
		11'd1234: begin
			vns_clockdomainsrenamer1_liteethudp_sel <= 1'd1;
		end
		default: begin
			vns_clockdomainsrenamer1_liteethudp_sel <= 1'd0;
		end
	endcase
end
assign soc_videooverlaysoc_packet_tx_cdc_asyncfifo_din = {soc_videooverlaysoc_packet_tx_cdc_fifo_in_last, soc_videooverlaysoc_packet_tx_cdc_fifo_in_first, soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_length, soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_ip_address, soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_dst_port, soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_src_port, soc_videooverlaysoc_packet_tx_cdc_fifo_in_payload_error, soc_videooverlaysoc_packet_tx_cdc_fifo_in_payload_data};
assign {soc_videooverlaysoc_packet_tx_cdc_fifo_out_last, soc_videooverlaysoc_packet_tx_cdc_fifo_out_first, soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_length, soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_ip_address, soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_dst_port, soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_src_port, soc_videooverlaysoc_packet_tx_cdc_fifo_out_payload_error, soc_videooverlaysoc_packet_tx_cdc_fifo_out_payload_data} = soc_videooverlaysoc_packet_tx_cdc_asyncfifo_dout;
assign soc_videooverlaysoc_packet_tx_cdc_sink_ready = soc_videooverlaysoc_packet_tx_cdc_asyncfifo_writable;
assign soc_videooverlaysoc_packet_tx_cdc_asyncfifo_we = soc_videooverlaysoc_packet_tx_cdc_sink_valid;
assign soc_videooverlaysoc_packet_tx_cdc_fifo_in_first = soc_videooverlaysoc_packet_tx_cdc_sink_first;
assign soc_videooverlaysoc_packet_tx_cdc_fifo_in_last = soc_videooverlaysoc_packet_tx_cdc_sink_last;
assign soc_videooverlaysoc_packet_tx_cdc_fifo_in_payload_data = soc_videooverlaysoc_packet_tx_cdc_sink_payload_data;
assign soc_videooverlaysoc_packet_tx_cdc_fifo_in_payload_error = soc_videooverlaysoc_packet_tx_cdc_sink_payload_error;
assign soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_src_port = soc_videooverlaysoc_packet_tx_cdc_sink_param_src_port;
assign soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_dst_port = soc_videooverlaysoc_packet_tx_cdc_sink_param_dst_port;
assign soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_ip_address = soc_videooverlaysoc_packet_tx_cdc_sink_param_ip_address;
assign soc_videooverlaysoc_packet_tx_cdc_fifo_in_param_length = soc_videooverlaysoc_packet_tx_cdc_sink_param_length;
assign soc_videooverlaysoc_packet_tx_cdc_source_valid = soc_videooverlaysoc_packet_tx_cdc_asyncfifo_readable;
assign soc_videooverlaysoc_packet_tx_cdc_source_first = soc_videooverlaysoc_packet_tx_cdc_fifo_out_first;
assign soc_videooverlaysoc_packet_tx_cdc_source_last = soc_videooverlaysoc_packet_tx_cdc_fifo_out_last;
assign soc_videooverlaysoc_packet_tx_cdc_source_payload_data = soc_videooverlaysoc_packet_tx_cdc_fifo_out_payload_data;
assign soc_videooverlaysoc_packet_tx_cdc_source_payload_error = soc_videooverlaysoc_packet_tx_cdc_fifo_out_payload_error;
assign soc_videooverlaysoc_packet_tx_cdc_source_param_src_port = soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_src_port;
assign soc_videooverlaysoc_packet_tx_cdc_source_param_dst_port = soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_dst_port;
assign soc_videooverlaysoc_packet_tx_cdc_source_param_ip_address = soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_ip_address;
assign soc_videooverlaysoc_packet_tx_cdc_source_param_length = soc_videooverlaysoc_packet_tx_cdc_fifo_out_param_length;
assign soc_videooverlaysoc_packet_tx_cdc_asyncfifo_re = soc_videooverlaysoc_packet_tx_cdc_source_ready;
assign soc_videooverlaysoc_packet_tx_cdc_graycounter0_ce = (soc_videooverlaysoc_packet_tx_cdc_asyncfifo_writable & soc_videooverlaysoc_packet_tx_cdc_asyncfifo_we);
assign soc_videooverlaysoc_packet_tx_cdc_graycounter1_ce = (soc_videooverlaysoc_packet_tx_cdc_asyncfifo_readable & soc_videooverlaysoc_packet_tx_cdc_asyncfifo_re);
assign soc_videooverlaysoc_packet_tx_cdc_asyncfifo_writable = (((soc_videooverlaysoc_packet_tx_cdc_graycounter0_q[2] == soc_videooverlaysoc_packet_tx_cdc_consume_wdomain[2]) | (soc_videooverlaysoc_packet_tx_cdc_graycounter0_q[1] == soc_videooverlaysoc_packet_tx_cdc_consume_wdomain[1])) | (soc_videooverlaysoc_packet_tx_cdc_graycounter0_q[0] != soc_videooverlaysoc_packet_tx_cdc_consume_wdomain[0]));
assign soc_videooverlaysoc_packet_tx_cdc_asyncfifo_readable = (soc_videooverlaysoc_packet_tx_cdc_graycounter1_q != soc_videooverlaysoc_packet_tx_cdc_produce_rdomain);
assign soc_videooverlaysoc_packet_tx_cdc_wrport_adr = soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_binary[1:0];
assign soc_videooverlaysoc_packet_tx_cdc_wrport_dat_w = soc_videooverlaysoc_packet_tx_cdc_asyncfifo_din;
assign soc_videooverlaysoc_packet_tx_cdc_wrport_we = soc_videooverlaysoc_packet_tx_cdc_graycounter0_ce;
assign soc_videooverlaysoc_packet_tx_cdc_rdport_adr = soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next_binary[1:0];
assign soc_videooverlaysoc_packet_tx_cdc_asyncfifo_dout = soc_videooverlaysoc_packet_tx_cdc_rdport_dat_r;
always @(*) begin
	soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_next_binary <= 3'd0;
	if (soc_videooverlaysoc_packet_tx_cdc_graycounter0_ce) begin
		soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_next_binary <= (soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_next_binary <= soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_binary;
	end
end
assign soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_next = (soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_next_binary ^ soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_next_binary[2:1]);
always @(*) begin
	soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next_binary <= 3'd0;
	if (soc_videooverlaysoc_packet_tx_cdc_graycounter1_ce) begin
		soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next_binary <= (soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next_binary <= soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_binary;
	end
end
assign soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next = (soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next_binary ^ soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next_binary[2:1]);
assign soc_videooverlaysoc_packet_tx_converter_converter_sink_valid = soc_videooverlaysoc_packet_tx_converter_sink_valid;
assign soc_videooverlaysoc_packet_tx_converter_converter_sink_first = soc_videooverlaysoc_packet_tx_converter_sink_first;
assign soc_videooverlaysoc_packet_tx_converter_converter_sink_last = soc_videooverlaysoc_packet_tx_converter_sink_last;
assign soc_videooverlaysoc_packet_tx_converter_sink_ready = soc_videooverlaysoc_packet_tx_converter_converter_sink_ready;
always @(*) begin
	soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data <= 36'd0;
	soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[7:0] <= soc_videooverlaysoc_packet_tx_converter_sink_payload_data[7:0];
	soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[8] <= soc_videooverlaysoc_packet_tx_converter_sink_payload_error[0];
	soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[16:9] <= soc_videooverlaysoc_packet_tx_converter_sink_payload_data[15:8];
	soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[17] <= soc_videooverlaysoc_packet_tx_converter_sink_payload_error[1];
	soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[25:18] <= soc_videooverlaysoc_packet_tx_converter_sink_payload_data[23:16];
	soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[26] <= soc_videooverlaysoc_packet_tx_converter_sink_payload_error[2];
	soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[34:27] <= soc_videooverlaysoc_packet_tx_converter_sink_payload_data[31:24];
	soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[35] <= soc_videooverlaysoc_packet_tx_converter_sink_payload_error[3];
end
assign soc_videooverlaysoc_packet_tx_converter_source_valid = soc_videooverlaysoc_packet_tx_converter_source_source_valid;
assign soc_videooverlaysoc_packet_tx_converter_source_first = soc_videooverlaysoc_packet_tx_converter_source_source_first;
assign soc_videooverlaysoc_packet_tx_converter_source_last = soc_videooverlaysoc_packet_tx_converter_source_source_last;
assign soc_videooverlaysoc_packet_tx_converter_source_source_ready = soc_videooverlaysoc_packet_tx_converter_source_ready;
assign {soc_videooverlaysoc_packet_tx_converter_source_payload_error, soc_videooverlaysoc_packet_tx_converter_source_payload_data} = soc_videooverlaysoc_packet_tx_converter_source_source_payload_data;
assign soc_videooverlaysoc_packet_tx_converter_source_param_src_port = soc_videooverlaysoc_packet_tx_converter_sink_param_src_port;
assign soc_videooverlaysoc_packet_tx_converter_source_param_dst_port = soc_videooverlaysoc_packet_tx_converter_sink_param_dst_port;
assign soc_videooverlaysoc_packet_tx_converter_source_param_ip_address = soc_videooverlaysoc_packet_tx_converter_sink_param_ip_address;
assign soc_videooverlaysoc_packet_tx_converter_source_param_length = soc_videooverlaysoc_packet_tx_converter_sink_param_length;
assign soc_videooverlaysoc_packet_tx_converter_source_source_valid = soc_videooverlaysoc_packet_tx_converter_converter_source_valid;
assign soc_videooverlaysoc_packet_tx_converter_converter_source_ready = soc_videooverlaysoc_packet_tx_converter_source_source_ready;
assign soc_videooverlaysoc_packet_tx_converter_source_source_first = soc_videooverlaysoc_packet_tx_converter_converter_source_first;
assign soc_videooverlaysoc_packet_tx_converter_source_source_last = soc_videooverlaysoc_packet_tx_converter_converter_source_last;
assign soc_videooverlaysoc_packet_tx_converter_source_source_payload_data = soc_videooverlaysoc_packet_tx_converter_converter_source_payload_data;
assign soc_videooverlaysoc_packet_tx_converter_converter_first = (soc_videooverlaysoc_packet_tx_converter_converter_mux == 1'd0);
assign soc_videooverlaysoc_packet_tx_converter_converter_last = (soc_videooverlaysoc_packet_tx_converter_converter_mux == 2'd3);
assign soc_videooverlaysoc_packet_tx_converter_converter_source_valid = soc_videooverlaysoc_packet_tx_converter_converter_sink_valid;
assign soc_videooverlaysoc_packet_tx_converter_converter_source_first = (soc_videooverlaysoc_packet_tx_converter_converter_sink_first & soc_videooverlaysoc_packet_tx_converter_converter_first);
assign soc_videooverlaysoc_packet_tx_converter_converter_source_last = (soc_videooverlaysoc_packet_tx_converter_converter_sink_last & soc_videooverlaysoc_packet_tx_converter_converter_last);
assign soc_videooverlaysoc_packet_tx_converter_converter_sink_ready = (soc_videooverlaysoc_packet_tx_converter_converter_last & soc_videooverlaysoc_packet_tx_converter_converter_source_ready);
always @(*) begin
	soc_videooverlaysoc_packet_tx_converter_converter_source_payload_data <= 9'd0;
	case (soc_videooverlaysoc_packet_tx_converter_converter_mux)
		1'd0: begin
			soc_videooverlaysoc_packet_tx_converter_converter_source_payload_data <= soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[8:0];
		end
		1'd1: begin
			soc_videooverlaysoc_packet_tx_converter_converter_source_payload_data <= soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[17:9];
		end
		2'd2: begin
			soc_videooverlaysoc_packet_tx_converter_converter_source_payload_data <= soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[26:18];
		end
		default: begin
			soc_videooverlaysoc_packet_tx_converter_converter_source_payload_data <= soc_videooverlaysoc_packet_tx_converter_converter_sink_payload_data[35:27];
		end
	endcase
end
assign soc_videooverlaysoc_packet_tx_converter_converter_source_payload_valid_token_count = soc_videooverlaysoc_packet_tx_converter_converter_last;
assign soc_videooverlaysoc_packet_rx_converter_converter_sink_valid = soc_videooverlaysoc_packet_rx_converter_sink_valid;
assign soc_videooverlaysoc_packet_rx_converter_converter_sink_first = soc_videooverlaysoc_packet_rx_converter_sink_first;
assign soc_videooverlaysoc_packet_rx_converter_converter_sink_last = soc_videooverlaysoc_packet_rx_converter_sink_last;
assign soc_videooverlaysoc_packet_rx_converter_sink_ready = soc_videooverlaysoc_packet_rx_converter_converter_sink_ready;
assign soc_videooverlaysoc_packet_rx_converter_converter_sink_payload_data = {soc_videooverlaysoc_packet_rx_converter_sink_payload_error, soc_videooverlaysoc_packet_rx_converter_sink_payload_data};
assign soc_videooverlaysoc_packet_rx_converter_source_valid = soc_videooverlaysoc_packet_rx_converter_source_source_valid;
assign soc_videooverlaysoc_packet_rx_converter_source_first = soc_videooverlaysoc_packet_rx_converter_source_source_first;
assign soc_videooverlaysoc_packet_rx_converter_source_last = soc_videooverlaysoc_packet_rx_converter_source_source_last;
assign soc_videooverlaysoc_packet_rx_converter_source_source_ready = soc_videooverlaysoc_packet_rx_converter_source_ready;
always @(*) begin
	soc_videooverlaysoc_packet_rx_converter_source_payload_data <= 32'd0;
	soc_videooverlaysoc_packet_rx_converter_source_payload_data[7:0] <= soc_videooverlaysoc_packet_rx_converter_source_source_payload_data[7:0];
	soc_videooverlaysoc_packet_rx_converter_source_payload_data[15:8] <= soc_videooverlaysoc_packet_rx_converter_source_source_payload_data[16:9];
	soc_videooverlaysoc_packet_rx_converter_source_payload_data[23:16] <= soc_videooverlaysoc_packet_rx_converter_source_source_payload_data[25:18];
	soc_videooverlaysoc_packet_rx_converter_source_payload_data[31:24] <= soc_videooverlaysoc_packet_rx_converter_source_source_payload_data[34:27];
end
always @(*) begin
	soc_videooverlaysoc_packet_rx_converter_source_payload_error <= 4'd0;
	soc_videooverlaysoc_packet_rx_converter_source_payload_error[0] <= soc_videooverlaysoc_packet_rx_converter_source_source_payload_data[8];
	soc_videooverlaysoc_packet_rx_converter_source_payload_error[1] <= soc_videooverlaysoc_packet_rx_converter_source_source_payload_data[17];
	soc_videooverlaysoc_packet_rx_converter_source_payload_error[2] <= soc_videooverlaysoc_packet_rx_converter_source_source_payload_data[26];
	soc_videooverlaysoc_packet_rx_converter_source_payload_error[3] <= soc_videooverlaysoc_packet_rx_converter_source_source_payload_data[35];
end
assign soc_videooverlaysoc_packet_rx_converter_source_source_valid = soc_videooverlaysoc_packet_rx_converter_converter_source_valid;
assign soc_videooverlaysoc_packet_rx_converter_converter_source_ready = soc_videooverlaysoc_packet_rx_converter_source_source_ready;
assign soc_videooverlaysoc_packet_rx_converter_source_source_first = soc_videooverlaysoc_packet_rx_converter_converter_source_first;
assign soc_videooverlaysoc_packet_rx_converter_source_source_last = soc_videooverlaysoc_packet_rx_converter_converter_source_last;
assign soc_videooverlaysoc_packet_rx_converter_source_source_payload_data = soc_videooverlaysoc_packet_rx_converter_converter_source_payload_data;
assign soc_videooverlaysoc_packet_rx_converter_converter_sink_ready = ((~soc_videooverlaysoc_packet_rx_converter_converter_strobe_all) | soc_videooverlaysoc_packet_rx_converter_converter_source_ready);
assign soc_videooverlaysoc_packet_rx_converter_converter_source_valid = soc_videooverlaysoc_packet_rx_converter_converter_strobe_all;
assign soc_videooverlaysoc_packet_rx_converter_converter_load_part = (soc_videooverlaysoc_packet_rx_converter_converter_sink_valid & soc_videooverlaysoc_packet_rx_converter_converter_sink_ready);
assign soc_videooverlaysoc_packet_rx_cdc_asyncfifo_din = {soc_videooverlaysoc_packet_rx_cdc_fifo_in_last, soc_videooverlaysoc_packet_rx_cdc_fifo_in_first, soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_length, soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_ip_address, soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_dst_port, soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_src_port, soc_videooverlaysoc_packet_rx_cdc_fifo_in_payload_error, soc_videooverlaysoc_packet_rx_cdc_fifo_in_payload_data};
assign {soc_videooverlaysoc_packet_rx_cdc_fifo_out_last, soc_videooverlaysoc_packet_rx_cdc_fifo_out_first, soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_length, soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_ip_address, soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_dst_port, soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_src_port, soc_videooverlaysoc_packet_rx_cdc_fifo_out_payload_error, soc_videooverlaysoc_packet_rx_cdc_fifo_out_payload_data} = soc_videooverlaysoc_packet_rx_cdc_asyncfifo_dout;
assign soc_videooverlaysoc_packet_rx_cdc_sink_ready = soc_videooverlaysoc_packet_rx_cdc_asyncfifo_writable;
assign soc_videooverlaysoc_packet_rx_cdc_asyncfifo_we = soc_videooverlaysoc_packet_rx_cdc_sink_valid;
assign soc_videooverlaysoc_packet_rx_cdc_fifo_in_first = soc_videooverlaysoc_packet_rx_cdc_sink_first;
assign soc_videooverlaysoc_packet_rx_cdc_fifo_in_last = soc_videooverlaysoc_packet_rx_cdc_sink_last;
assign soc_videooverlaysoc_packet_rx_cdc_fifo_in_payload_data = soc_videooverlaysoc_packet_rx_cdc_sink_payload_data;
assign soc_videooverlaysoc_packet_rx_cdc_fifo_in_payload_error = soc_videooverlaysoc_packet_rx_cdc_sink_payload_error;
assign soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_src_port = soc_videooverlaysoc_packet_rx_cdc_sink_param_src_port;
assign soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_dst_port = soc_videooverlaysoc_packet_rx_cdc_sink_param_dst_port;
assign soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_ip_address = soc_videooverlaysoc_packet_rx_cdc_sink_param_ip_address;
assign soc_videooverlaysoc_packet_rx_cdc_fifo_in_param_length = soc_videooverlaysoc_packet_rx_cdc_sink_param_length;
assign soc_videooverlaysoc_packet_rx_cdc_source_valid = soc_videooverlaysoc_packet_rx_cdc_asyncfifo_readable;
assign soc_videooverlaysoc_packet_rx_cdc_source_first = soc_videooverlaysoc_packet_rx_cdc_fifo_out_first;
assign soc_videooverlaysoc_packet_rx_cdc_source_last = soc_videooverlaysoc_packet_rx_cdc_fifo_out_last;
assign soc_videooverlaysoc_packet_rx_cdc_source_payload_data = soc_videooverlaysoc_packet_rx_cdc_fifo_out_payload_data;
assign soc_videooverlaysoc_packet_rx_cdc_source_payload_error = soc_videooverlaysoc_packet_rx_cdc_fifo_out_payload_error;
assign soc_videooverlaysoc_packet_rx_cdc_source_param_src_port = soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_src_port;
assign soc_videooverlaysoc_packet_rx_cdc_source_param_dst_port = soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_dst_port;
assign soc_videooverlaysoc_packet_rx_cdc_source_param_ip_address = soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_ip_address;
assign soc_videooverlaysoc_packet_rx_cdc_source_param_length = soc_videooverlaysoc_packet_rx_cdc_fifo_out_param_length;
assign soc_videooverlaysoc_packet_rx_cdc_asyncfifo_re = soc_videooverlaysoc_packet_rx_cdc_source_ready;
assign soc_videooverlaysoc_packet_rx_cdc_graycounter0_ce = (soc_videooverlaysoc_packet_rx_cdc_asyncfifo_writable & soc_videooverlaysoc_packet_rx_cdc_asyncfifo_we);
assign soc_videooverlaysoc_packet_rx_cdc_graycounter1_ce = (soc_videooverlaysoc_packet_rx_cdc_asyncfifo_readable & soc_videooverlaysoc_packet_rx_cdc_asyncfifo_re);
assign soc_videooverlaysoc_packet_rx_cdc_asyncfifo_writable = (((soc_videooverlaysoc_packet_rx_cdc_graycounter0_q[2] == soc_videooverlaysoc_packet_rx_cdc_consume_wdomain[2]) | (soc_videooverlaysoc_packet_rx_cdc_graycounter0_q[1] == soc_videooverlaysoc_packet_rx_cdc_consume_wdomain[1])) | (soc_videooverlaysoc_packet_rx_cdc_graycounter0_q[0] != soc_videooverlaysoc_packet_rx_cdc_consume_wdomain[0]));
assign soc_videooverlaysoc_packet_rx_cdc_asyncfifo_readable = (soc_videooverlaysoc_packet_rx_cdc_graycounter1_q != soc_videooverlaysoc_packet_rx_cdc_produce_rdomain);
assign soc_videooverlaysoc_packet_rx_cdc_wrport_adr = soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_binary[1:0];
assign soc_videooverlaysoc_packet_rx_cdc_wrport_dat_w = soc_videooverlaysoc_packet_rx_cdc_asyncfifo_din;
assign soc_videooverlaysoc_packet_rx_cdc_wrport_we = soc_videooverlaysoc_packet_rx_cdc_graycounter0_ce;
assign soc_videooverlaysoc_packet_rx_cdc_rdport_adr = soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next_binary[1:0];
assign soc_videooverlaysoc_packet_rx_cdc_asyncfifo_dout = soc_videooverlaysoc_packet_rx_cdc_rdport_dat_r;
always @(*) begin
	soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_next_binary <= 3'd0;
	if (soc_videooverlaysoc_packet_rx_cdc_graycounter0_ce) begin
		soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_next_binary <= (soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_next_binary <= soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_binary;
	end
end
assign soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_next = (soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_next_binary ^ soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_next_binary[2:1]);
always @(*) begin
	soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next_binary <= 3'd0;
	if (soc_videooverlaysoc_packet_rx_cdc_graycounter1_ce) begin
		soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next_binary <= (soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next_binary <= soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_binary;
	end
end
assign soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next = (soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next_binary ^ soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next_binary[2:1]);
assign soc_videooverlaysoc_core_crossbar_source_valid = soc_videooverlaysoc_packet_internal_port_sink_valid;
assign soc_videooverlaysoc_packet_internal_port_sink_ready = soc_videooverlaysoc_core_crossbar_source_ready;
assign soc_videooverlaysoc_core_crossbar_source_first = soc_videooverlaysoc_packet_internal_port_sink_first;
assign soc_videooverlaysoc_core_crossbar_source_last = soc_videooverlaysoc_packet_internal_port_sink_last;
assign soc_videooverlaysoc_core_crossbar_source_payload_data = soc_videooverlaysoc_packet_internal_port_sink_payload_data;
assign soc_videooverlaysoc_core_crossbar_source_payload_error = soc_videooverlaysoc_packet_internal_port_sink_payload_error;
assign soc_videooverlaysoc_core_crossbar_source_param_src_port = soc_videooverlaysoc_packet_internal_port_sink_param_src_port;
assign soc_videooverlaysoc_core_crossbar_source_param_dst_port = soc_videooverlaysoc_packet_internal_port_sink_param_dst_port;
assign soc_videooverlaysoc_core_crossbar_source_param_ip_address = soc_videooverlaysoc_packet_internal_port_sink_param_ip_address;
assign soc_videooverlaysoc_core_crossbar_source_param_length = soc_videooverlaysoc_packet_internal_port_sink_param_length;
assign soc_videooverlaysoc_packet_internal_port_source_valid = soc_videooverlaysoc_core_crossbar_sink_valid;
assign soc_videooverlaysoc_core_crossbar_sink_ready = soc_videooverlaysoc_packet_internal_port_source_ready;
assign soc_videooverlaysoc_packet_internal_port_source_first = soc_videooverlaysoc_core_crossbar_sink_first;
assign soc_videooverlaysoc_packet_internal_port_source_last = soc_videooverlaysoc_core_crossbar_sink_last;
assign soc_videooverlaysoc_packet_internal_port_source_payload_data = soc_videooverlaysoc_core_crossbar_sink_payload_data;
assign soc_videooverlaysoc_packet_internal_port_source_payload_error = soc_videooverlaysoc_core_crossbar_sink_payload_error;
assign soc_videooverlaysoc_packet_internal_port_source_param_src_port = soc_videooverlaysoc_core_crossbar_sink_param_src_port;
assign soc_videooverlaysoc_packet_internal_port_source_param_dst_port = soc_videooverlaysoc_core_crossbar_sink_param_dst_port;
assign soc_videooverlaysoc_packet_internal_port_source_param_ip_address = soc_videooverlaysoc_core_crossbar_sink_param_ip_address;
assign soc_videooverlaysoc_packet_internal_port_source_param_length = soc_videooverlaysoc_core_crossbar_sink_param_length;
assign soc_videooverlaysoc_dispatcher_sel0 = (~soc_videooverlaysoc_packet_source_source_param_pf);
assign soc_videooverlaysoc_wishbone_sink_valid = soc_videooverlaysoc_record_receiver_source_source_valid;
assign soc_videooverlaysoc_record_receiver_source_source_ready = soc_videooverlaysoc_wishbone_sink_ready;
assign soc_videooverlaysoc_wishbone_sink_first = soc_videooverlaysoc_record_receiver_source_source_first;
assign soc_videooverlaysoc_wishbone_sink_last = soc_videooverlaysoc_record_receiver_source_source_last;
assign soc_videooverlaysoc_wishbone_sink_payload_addr = soc_videooverlaysoc_record_receiver_source_source_payload_addr;
assign soc_videooverlaysoc_wishbone_sink_payload_data = soc_videooverlaysoc_record_receiver_source_source_payload_data;
assign soc_videooverlaysoc_wishbone_sink_param_we = soc_videooverlaysoc_record_receiver_source_source_param_we;
assign soc_videooverlaysoc_wishbone_sink_param_count = soc_videooverlaysoc_record_receiver_source_source_param_count;
assign soc_videooverlaysoc_wishbone_sink_param_base_addr = soc_videooverlaysoc_record_receiver_source_source_param_base_addr;
assign soc_videooverlaysoc_wishbone_sink_param_be = soc_videooverlaysoc_record_receiver_source_source_param_be;
assign soc_videooverlaysoc_record_sender_sink_sink_valid = soc_videooverlaysoc_wishbone_source_valid;
assign soc_videooverlaysoc_wishbone_source_ready = soc_videooverlaysoc_record_sender_sink_sink_ready;
assign soc_videooverlaysoc_record_sender_sink_sink_first = soc_videooverlaysoc_wishbone_source_first;
assign soc_videooverlaysoc_record_sender_sink_sink_last = soc_videooverlaysoc_wishbone_source_last;
assign soc_videooverlaysoc_record_sender_sink_sink_payload_addr = soc_videooverlaysoc_wishbone_source_payload_addr;
assign soc_videooverlaysoc_record_sender_sink_sink_payload_data = soc_videooverlaysoc_wishbone_source_payload_data;
assign soc_videooverlaysoc_record_sender_sink_sink_param_we = soc_videooverlaysoc_wishbone_source_param_we;
assign soc_videooverlaysoc_record_sender_sink_sink_param_count = soc_videooverlaysoc_wishbone_source_param_count;
assign soc_videooverlaysoc_record_sender_sink_sink_param_base_addr = soc_videooverlaysoc_wishbone_source_param_base_addr;
assign soc_videooverlaysoc_record_sender_sink_sink_param_be = soc_videooverlaysoc_wishbone_source_param_be;
assign soc_videooverlaysoc_packet_user_port_sink_valid = soc_videooverlaysoc_packet_source_valid;
assign soc_videooverlaysoc_packet_source_ready = soc_videooverlaysoc_packet_user_port_sink_ready;
assign soc_videooverlaysoc_packet_user_port_sink_first = soc_videooverlaysoc_packet_source_first;
assign soc_videooverlaysoc_packet_user_port_sink_last = soc_videooverlaysoc_packet_source_last;
assign soc_videooverlaysoc_packet_user_port_sink_payload_data = soc_videooverlaysoc_packet_source_payload_data;
assign soc_videooverlaysoc_packet_user_port_sink_payload_error = soc_videooverlaysoc_packet_source_payload_error;
assign soc_videooverlaysoc_packet_user_port_sink_param_src_port = soc_videooverlaysoc_packet_source_param_src_port;
assign soc_videooverlaysoc_packet_user_port_sink_param_dst_port = soc_videooverlaysoc_packet_source_param_dst_port;
assign soc_videooverlaysoc_packet_user_port_sink_param_ip_address = soc_videooverlaysoc_packet_source_param_ip_address;
assign soc_videooverlaysoc_packet_user_port_sink_param_length = soc_videooverlaysoc_packet_source_param_length;
assign soc_videooverlaysoc_packet_sink_sink_valid = soc_videooverlaysoc_packet_user_port_source_valid;
assign soc_videooverlaysoc_packet_user_port_source_ready = soc_videooverlaysoc_packet_sink_sink_ready;
assign soc_videooverlaysoc_packet_sink_sink_first = soc_videooverlaysoc_packet_user_port_source_first;
assign soc_videooverlaysoc_packet_sink_sink_last = soc_videooverlaysoc_packet_user_port_source_last;
assign soc_videooverlaysoc_packet_sink_sink_payload_data = soc_videooverlaysoc_packet_user_port_source_payload_data;
assign soc_videooverlaysoc_packet_sink_sink_payload_error = soc_videooverlaysoc_packet_user_port_source_payload_error;
assign soc_videooverlaysoc_packet_sink_sink_param_src_port = soc_videooverlaysoc_packet_user_port_source_param_src_port;
assign soc_videooverlaysoc_packet_sink_sink_param_dst_port = soc_videooverlaysoc_packet_user_port_source_param_dst_port;
assign soc_videooverlaysoc_packet_sink_sink_param_ip_address = soc_videooverlaysoc_packet_user_port_source_param_ip_address;
assign soc_videooverlaysoc_packet_sink_sink_param_length = soc_videooverlaysoc_packet_user_port_source_param_length;
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_valid = soc_videooverlaysoc_packet_sink_valid;
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_last = soc_videooverlaysoc_packet_sink_last;
assign soc_videooverlaysoc_packet_sink_ready = soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_ready;
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_magic = 15'd20079;
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_port_size = 3'd4;
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_addr_size = 3'd4;
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_pf = soc_videooverlaysoc_packet_sink_param_pf;
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_pr = soc_videooverlaysoc_packet_sink_param_pr;
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_nr = soc_videooverlaysoc_packet_sink_param_nr;
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_version = 1'd1;
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_payload_data = soc_videooverlaysoc_packet_sink_payload_data;
always @(*) begin
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header <= 64'd0;
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header[31:28] <= {soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_addr_size[3:0]};
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header[15:0] <= {soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_magic[7:0], soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_magic[15:8]};
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header[18] <= {soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_nr};
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header[16] <= {soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_pf};
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header[27:24] <= {soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_port_size[3:0]};
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header[17] <= {soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_pr};
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header[23:20] <= {soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_param_version[3:0]};
end
assign soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_payload_error = soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_payload_error;
always @(*) begin
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_valid <= 1'd0;
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter_ce <= 1'd0;
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_last <= 1'd0;
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_payload_data <= 32'd0;
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_load <= 1'd0;
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_shift <= 1'd0;
	vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_next_state <= 2'd0;
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter_reset <= 1'd0;
	vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_next_state <= vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_state;
	case (vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_valid <= 1'd1;
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_last <= 1'd0;
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_payload_data <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header_reg[63:32];
			if ((soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_valid & soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_ready)) begin
				soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_shift <= 1'd1;
				soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter_ce <= 1'd1;
				if ((soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter == 1'd0)) begin
					vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_valid <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_valid;
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_last <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_last;
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_payload_data <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_payload_data;
			if ((soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_valid & soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_ready)) begin
				soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_ready <= 1'd1;
				if (soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_last) begin
					vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_valid) begin
				soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_sink_ready <= 1'd0;
				soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_valid <= 1'd1;
				soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_last <= 1'd0;
				soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_payload_data <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header[31:0];
				if ((soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_valid & soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_ready)) begin
					soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_load <= 1'd1;
					vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_next_state <= 1'd1;
				end
			end
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_packet_source_param_dst_port <= 16'd0;
	soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_ready <= 1'd0;
	soc_videooverlaysoc_packet_source_param_ip_address <= 32'd0;
	soc_videooverlaysoc_packet_source_param_length <= 16'd0;
	vns_liteethetherbonepackettx_fsm_next_state <= 1'd0;
	soc_videooverlaysoc_packet_source_valid <= 1'd0;
	soc_videooverlaysoc_packet_source_first <= 1'd0;
	soc_videooverlaysoc_packet_source_last <= 1'd0;
	soc_videooverlaysoc_packet_source_payload_data <= 32'd0;
	soc_videooverlaysoc_packet_source_payload_error <= 4'd0;
	soc_videooverlaysoc_packet_source_param_src_port <= 16'd0;
	vns_liteethetherbonepackettx_fsm_next_state <= vns_liteethetherbonepackettx_fsm_state;
	case (vns_liteethetherbonepackettx_fsm_state)
		1'd1: begin
			soc_videooverlaysoc_packet_source_valid <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_valid;
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_ready <= soc_videooverlaysoc_packet_source_ready;
			soc_videooverlaysoc_packet_source_first <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_first;
			soc_videooverlaysoc_packet_source_last <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_last;
			soc_videooverlaysoc_packet_source_payload_data <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_payload_data;
			soc_videooverlaysoc_packet_source_payload_error <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_payload_error;
			soc_videooverlaysoc_packet_source_param_src_port <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_param_src_port;
			soc_videooverlaysoc_packet_source_param_dst_port <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_param_dst_port;
			soc_videooverlaysoc_packet_source_param_ip_address <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_param_ip_address;
			soc_videooverlaysoc_packet_source_param_length <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_param_length;
			soc_videooverlaysoc_packet_source_param_src_port <= 11'd1234;
			soc_videooverlaysoc_packet_source_param_dst_port <= 11'd1234;
			soc_videooverlaysoc_packet_source_param_ip_address <= soc_videooverlaysoc_packet_sink_param_ip_address;
			soc_videooverlaysoc_packet_source_param_length <= (soc_videooverlaysoc_packet_sink_param_length + 4'd8);
			if (((soc_videooverlaysoc_packet_source_valid & soc_videooverlaysoc_packet_source_last) & soc_videooverlaysoc_packet_source_ready)) begin
				vns_liteethetherbonepackettx_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_ready <= 1'd1;
			if (soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_valid) begin
				soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_source_ready <= 1'd0;
				vns_liteethetherbonepackettx_fsm_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_packet_depacketizer_sink_valid = soc_videooverlaysoc_packet_sink_sink_valid;
assign soc_videooverlaysoc_packet_sink_sink_ready = soc_videooverlaysoc_packet_depacketizer_sink_ready;
assign soc_videooverlaysoc_packet_depacketizer_sink_first = soc_videooverlaysoc_packet_sink_sink_first;
assign soc_videooverlaysoc_packet_depacketizer_sink_last = soc_videooverlaysoc_packet_sink_sink_last;
assign soc_videooverlaysoc_packet_depacketizer_sink_payload_data = soc_videooverlaysoc_packet_sink_sink_payload_data;
assign soc_videooverlaysoc_packet_depacketizer_sink_payload_error = soc_videooverlaysoc_packet_sink_sink_payload_error;
assign soc_videooverlaysoc_packet_depacketizer_sink_param_src_port = soc_videooverlaysoc_packet_sink_sink_param_src_port;
assign soc_videooverlaysoc_packet_depacketizer_sink_param_dst_port = soc_videooverlaysoc_packet_sink_sink_param_dst_port;
assign soc_videooverlaysoc_packet_depacketizer_sink_param_ip_address = soc_videooverlaysoc_packet_sink_sink_param_ip_address;
assign soc_videooverlaysoc_packet_depacketizer_sink_param_length = soc_videooverlaysoc_packet_sink_sink_param_length;
assign soc_videooverlaysoc_packet_source_source_last = soc_videooverlaysoc_packet_depacketizer_source_last;
assign soc_videooverlaysoc_packet_source_source_param_pf = soc_videooverlaysoc_packet_depacketizer_source_param_pf;
assign soc_videooverlaysoc_packet_source_source_param_pr = soc_videooverlaysoc_packet_depacketizer_source_param_pr;
assign soc_videooverlaysoc_packet_source_source_param_nr = soc_videooverlaysoc_packet_depacketizer_source_param_nr;
assign soc_videooverlaysoc_packet_source_source_payload_data = soc_videooverlaysoc_packet_depacketizer_source_payload_data;
assign soc_videooverlaysoc_packet_source_source_param_src_port = soc_videooverlaysoc_packet_sink_sink_param_src_port;
assign soc_videooverlaysoc_packet_source_source_param_dst_port = soc_videooverlaysoc_packet_sink_sink_param_dst_port;
assign soc_videooverlaysoc_packet_source_source_param_ip_address = soc_videooverlaysoc_packet_sink_sink_param_ip_address;
assign soc_videooverlaysoc_packet_source_source_param_length = (soc_videooverlaysoc_packet_sink_sink_param_length - 4'd8);
assign soc_videooverlaysoc_packet_depacketizer_header = soc_videooverlaysoc_packet_depacketizer_header_reg;
assign soc_videooverlaysoc_packet_depacketizer_source_payload_error = soc_videooverlaysoc_packet_depacketizer_sink_payload_error;
assign soc_videooverlaysoc_packet_depacketizer_source_last = (soc_videooverlaysoc_packet_depacketizer_sink_last | soc_videooverlaysoc_packet_depacketizer_no_payload);
assign soc_videooverlaysoc_packet_depacketizer_source_payload_data = soc_videooverlaysoc_packet_depacketizer_sink_payload_data;
assign soc_videooverlaysoc_packet_depacketizer_source_param_addr_size = {vns_slice_proxy76[3:0]};
assign soc_videooverlaysoc_packet_depacketizer_source_param_magic = {vns_slice_proxy78[7:0], vns_slice_proxy77[15:8]};
assign soc_videooverlaysoc_packet_depacketizer_source_param_nr = {vns_slice_proxy79};
assign soc_videooverlaysoc_packet_depacketizer_source_param_pf = {vns_slice_proxy80};
assign soc_videooverlaysoc_packet_depacketizer_source_param_port_size = {vns_slice_proxy81[3:0]};
assign soc_videooverlaysoc_packet_depacketizer_source_param_pr = {vns_slice_proxy82};
assign soc_videooverlaysoc_packet_depacketizer_source_param_version = {vns_slice_proxy83[3:0]};
always @(*) begin
	soc_videooverlaysoc_packet_depacketizer_shift <= 1'd0;
	soc_videooverlaysoc_packet_depacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_packet_depacketizer_source_valid <= 1'd0;
	soc_videooverlaysoc_packet_depacketizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_packet_depacketizer_counter_ce <= 1'd0;
	vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_next_state <= 2'd0;
	vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_next_state <= vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_state;
	case (vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_packet_depacketizer_sink_ready <= 1'd1;
			if (soc_videooverlaysoc_packet_depacketizer_sink_valid) begin
				soc_videooverlaysoc_packet_depacketizer_counter_ce <= 1'd1;
				soc_videooverlaysoc_packet_depacketizer_shift <= 1'd1;
				if ((soc_videooverlaysoc_packet_depacketizer_counter == 1'd0)) begin
					vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_packet_depacketizer_sink_ready <= soc_videooverlaysoc_packet_depacketizer_source_ready;
			soc_videooverlaysoc_packet_depacketizer_source_valid <= (soc_videooverlaysoc_packet_depacketizer_sink_valid | soc_videooverlaysoc_packet_depacketizer_no_payload);
			if (((soc_videooverlaysoc_packet_depacketizer_source_valid & soc_videooverlaysoc_packet_depacketizer_source_ready) & soc_videooverlaysoc_packet_depacketizer_source_last)) begin
				vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_packet_depacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_packet_depacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_packet_depacketizer_sink_valid) begin
				soc_videooverlaysoc_packet_depacketizer_shift <= 1'd1;
				vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_packet_depacketizer_is_el = ((~(vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_state == 2'd2)) & (vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_next_state == 2'd2));
always @(*) begin
	soc_videooverlaysoc_packet_source_source_valid <= 1'd0;
	vns_liteethetherbonepacketrx_fsm_next_state <= 2'd0;
	soc_videooverlaysoc_packet_depacketizer_source_ready <= 1'd0;
	vns_liteethetherbonepacketrx_fsm_next_state <= vns_liteethetherbonepacketrx_fsm_state;
	case (vns_liteethetherbonepacketrx_fsm_state)
		1'd1: begin
			if (soc_videooverlaysoc_packet_valid) begin
				vns_liteethetherbonepacketrx_fsm_next_state <= 2'd2;
			end else begin
				vns_liteethetherbonepacketrx_fsm_next_state <= 2'd3;
			end
		end
		2'd2: begin
			soc_videooverlaysoc_packet_source_source_valid <= soc_videooverlaysoc_packet_depacketizer_source_valid;
			soc_videooverlaysoc_packet_depacketizer_source_ready <= soc_videooverlaysoc_packet_source_source_ready;
			if (((soc_videooverlaysoc_packet_source_source_valid & soc_videooverlaysoc_packet_source_source_last) & soc_videooverlaysoc_packet_source_source_ready)) begin
				vns_liteethetherbonepacketrx_fsm_next_state <= 1'd0;
			end
		end
		2'd3: begin
			soc_videooverlaysoc_packet_depacketizer_source_ready <= 1'd1;
			if (((soc_videooverlaysoc_packet_depacketizer_source_valid & soc_videooverlaysoc_packet_depacketizer_source_last) & soc_videooverlaysoc_packet_depacketizer_source_ready)) begin
				vns_liteethetherbonepacketrx_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_packet_depacketizer_source_ready <= 1'd1;
			if (soc_videooverlaysoc_packet_depacketizer_source_valid) begin
				soc_videooverlaysoc_packet_depacketizer_source_ready <= 1'd0;
				vns_liteethetherbonepacketrx_fsm_next_state <= 1'd1;
			end
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_probe_source_param_addr_size <= 4'd0;
	soc_videooverlaysoc_probe_source_param_nr <= 1'd0;
	soc_videooverlaysoc_probe_source_param_pf <= 1'd0;
	soc_videooverlaysoc_probe_source_param_port_size <= 4'd0;
	soc_videooverlaysoc_probe_source_param_pr <= 1'd0;
	vns_liteethetherboneprobe_next_state <= 1'd0;
	soc_videooverlaysoc_probe_source_param_src_port <= 16'd0;
	soc_videooverlaysoc_probe_source_param_dst_port <= 16'd0;
	soc_videooverlaysoc_probe_source_param_ip_address <= 32'd0;
	soc_videooverlaysoc_probe_source_param_length <= 16'd0;
	soc_videooverlaysoc_probe_sink_ready <= 1'd0;
	soc_videooverlaysoc_probe_source_valid <= 1'd0;
	soc_videooverlaysoc_probe_source_first <= 1'd0;
	soc_videooverlaysoc_probe_source_last <= 1'd0;
	soc_videooverlaysoc_probe_source_payload_data <= 32'd0;
	soc_videooverlaysoc_probe_source_payload_error <= 4'd0;
	vns_liteethetherboneprobe_next_state <= vns_liteethetherboneprobe_state;
	case (vns_liteethetherboneprobe_state)
		1'd1: begin
			soc_videooverlaysoc_probe_source_valid <= soc_videooverlaysoc_probe_sink_valid;
			soc_videooverlaysoc_probe_sink_ready <= soc_videooverlaysoc_probe_source_ready;
			soc_videooverlaysoc_probe_source_first <= soc_videooverlaysoc_probe_sink_first;
			soc_videooverlaysoc_probe_source_last <= soc_videooverlaysoc_probe_sink_last;
			soc_videooverlaysoc_probe_source_payload_data <= soc_videooverlaysoc_probe_sink_payload_data;
			soc_videooverlaysoc_probe_source_payload_error <= soc_videooverlaysoc_probe_sink_payload_error;
			soc_videooverlaysoc_probe_source_param_addr_size <= soc_videooverlaysoc_probe_sink_param_addr_size;
			soc_videooverlaysoc_probe_source_param_nr <= soc_videooverlaysoc_probe_sink_param_nr;
			soc_videooverlaysoc_probe_source_param_pf <= soc_videooverlaysoc_probe_sink_param_pf;
			soc_videooverlaysoc_probe_source_param_port_size <= soc_videooverlaysoc_probe_sink_param_port_size;
			soc_videooverlaysoc_probe_source_param_pr <= soc_videooverlaysoc_probe_sink_param_pr;
			soc_videooverlaysoc_probe_source_param_src_port <= soc_videooverlaysoc_probe_sink_param_src_port;
			soc_videooverlaysoc_probe_source_param_dst_port <= soc_videooverlaysoc_probe_sink_param_dst_port;
			soc_videooverlaysoc_probe_source_param_ip_address <= soc_videooverlaysoc_probe_sink_param_ip_address;
			soc_videooverlaysoc_probe_source_param_length <= soc_videooverlaysoc_probe_sink_param_length;
			soc_videooverlaysoc_probe_source_param_pf <= 1'd0;
			soc_videooverlaysoc_probe_source_param_pr <= 1'd1;
			if (((soc_videooverlaysoc_probe_source_valid & soc_videooverlaysoc_probe_source_last) & soc_videooverlaysoc_probe_source_ready)) begin
				vns_liteethetherboneprobe_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_probe_sink_ready <= 1'd1;
			if (soc_videooverlaysoc_probe_sink_valid) begin
				soc_videooverlaysoc_probe_sink_ready <= 1'd0;
				vns_liteethetherboneprobe_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_record_depacketizer_sink_valid = soc_videooverlaysoc_record_sink_sink_valid;
assign soc_videooverlaysoc_record_sink_sink_ready = soc_videooverlaysoc_record_depacketizer_sink_ready;
assign soc_videooverlaysoc_record_depacketizer_sink_first = soc_videooverlaysoc_record_sink_sink_first;
assign soc_videooverlaysoc_record_depacketizer_sink_last = soc_videooverlaysoc_record_sink_sink_last;
assign soc_videooverlaysoc_record_depacketizer_sink_payload_data = soc_videooverlaysoc_record_sink_sink_payload_data;
assign soc_videooverlaysoc_record_depacketizer_sink_payload_error = soc_videooverlaysoc_record_sink_sink_payload_error;
assign soc_videooverlaysoc_record_depacketizer_sink_param_addr_size = soc_videooverlaysoc_record_sink_sink_param_addr_size;
assign soc_videooverlaysoc_record_depacketizer_sink_param_nr = soc_videooverlaysoc_record_sink_sink_param_nr;
assign soc_videooverlaysoc_record_depacketizer_sink_param_pf = soc_videooverlaysoc_record_sink_sink_param_pf;
assign soc_videooverlaysoc_record_depacketizer_sink_param_port_size = soc_videooverlaysoc_record_sink_sink_param_port_size;
assign soc_videooverlaysoc_record_depacketizer_sink_param_pr = soc_videooverlaysoc_record_sink_sink_param_pr;
assign soc_videooverlaysoc_record_depacketizer_sink_param_src_port = soc_videooverlaysoc_record_sink_sink_param_src_port;
assign soc_videooverlaysoc_record_depacketizer_sink_param_dst_port = soc_videooverlaysoc_record_sink_sink_param_dst_port;
assign soc_videooverlaysoc_record_depacketizer_sink_param_ip_address = soc_videooverlaysoc_record_sink_sink_param_ip_address;
assign soc_videooverlaysoc_record_depacketizer_sink_param_length = soc_videooverlaysoc_record_sink_sink_param_length;
assign soc_videooverlaysoc_record_receiver_sink_sink_valid = soc_videooverlaysoc_record_depacketizer_source_valid;
assign soc_videooverlaysoc_record_depacketizer_source_ready = soc_videooverlaysoc_record_receiver_sink_sink_ready;
assign soc_videooverlaysoc_record_receiver_sink_sink_first = soc_videooverlaysoc_record_depacketizer_source_first;
assign soc_videooverlaysoc_record_receiver_sink_sink_last = soc_videooverlaysoc_record_depacketizer_source_last;
assign soc_videooverlaysoc_record_receiver_sink_sink_payload_error = soc_videooverlaysoc_record_depacketizer_source_payload_error;
assign soc_videooverlaysoc_record_receiver_sink_sink_param_bca = soc_videooverlaysoc_record_depacketizer_source_param_bca;
assign soc_videooverlaysoc_record_receiver_sink_sink_param_byte_enable = soc_videooverlaysoc_record_depacketizer_source_param_byte_enable;
assign soc_videooverlaysoc_record_receiver_sink_sink_param_cyc = soc_videooverlaysoc_record_depacketizer_source_param_cyc;
assign soc_videooverlaysoc_record_receiver_sink_sink_param_rca = soc_videooverlaysoc_record_depacketizer_source_param_rca;
assign soc_videooverlaysoc_record_receiver_sink_sink_param_rcount = soc_videooverlaysoc_record_depacketizer_source_param_rcount;
assign soc_videooverlaysoc_record_receiver_sink_sink_param_rff = soc_videooverlaysoc_record_depacketizer_source_param_rff;
assign soc_videooverlaysoc_record_receiver_sink_sink_param_wca = soc_videooverlaysoc_record_depacketizer_source_param_wca;
assign soc_videooverlaysoc_record_receiver_sink_sink_param_wcount = soc_videooverlaysoc_record_depacketizer_source_param_wcount;
assign soc_videooverlaysoc_record_receiver_sink_sink_param_wff = soc_videooverlaysoc_record_depacketizer_source_param_wff;
always @(*) begin
	soc_videooverlaysoc_record_receiver_sink_sink_payload_data <= 32'd0;
	soc_videooverlaysoc_record_receiver_sink_sink_payload_data <= soc_videooverlaysoc_record_depacketizer_source_payload_data;
	soc_videooverlaysoc_record_receiver_sink_sink_payload_data <= {soc_videooverlaysoc_record_depacketizer_source_payload_data[7:0], soc_videooverlaysoc_record_depacketizer_source_payload_data[15:8], soc_videooverlaysoc_record_depacketizer_source_payload_data[23:16], soc_videooverlaysoc_record_depacketizer_source_payload_data[31:24]};
end
assign soc_videooverlaysoc_record_packetizer_sink_valid = soc_videooverlaysoc_record_sender_source_source_valid;
assign soc_videooverlaysoc_record_sender_source_source_ready = soc_videooverlaysoc_record_packetizer_sink_ready;
assign soc_videooverlaysoc_record_packetizer_sink_first = soc_videooverlaysoc_record_sender_source_source_first;
assign soc_videooverlaysoc_record_packetizer_sink_last = soc_videooverlaysoc_record_sender_source_source_last;
assign soc_videooverlaysoc_record_packetizer_sink_payload_error = soc_videooverlaysoc_record_sender_source_source_payload_error;
assign soc_videooverlaysoc_record_packetizer_sink_param_bca = soc_videooverlaysoc_record_sender_source_source_param_bca;
assign soc_videooverlaysoc_record_packetizer_sink_param_byte_enable = soc_videooverlaysoc_record_sender_source_source_param_byte_enable;
assign soc_videooverlaysoc_record_packetizer_sink_param_cyc = soc_videooverlaysoc_record_sender_source_source_param_cyc;
assign soc_videooverlaysoc_record_packetizer_sink_param_rca = soc_videooverlaysoc_record_sender_source_source_param_rca;
assign soc_videooverlaysoc_record_packetizer_sink_param_rcount = soc_videooverlaysoc_record_sender_source_source_param_rcount;
assign soc_videooverlaysoc_record_packetizer_sink_param_rff = soc_videooverlaysoc_record_sender_source_source_param_rff;
assign soc_videooverlaysoc_record_packetizer_sink_param_wca = soc_videooverlaysoc_record_sender_source_source_param_wca;
assign soc_videooverlaysoc_record_packetizer_sink_param_wcount = soc_videooverlaysoc_record_sender_source_source_param_wcount;
assign soc_videooverlaysoc_record_packetizer_sink_param_wff = soc_videooverlaysoc_record_sender_source_source_param_wff;
assign soc_videooverlaysoc_record_source_source_valid = soc_videooverlaysoc_record_packetizer_source_valid;
assign soc_videooverlaysoc_record_packetizer_source_ready = soc_videooverlaysoc_record_source_source_ready;
assign soc_videooverlaysoc_record_source_source_first = soc_videooverlaysoc_record_packetizer_source_first;
assign soc_videooverlaysoc_record_source_source_last = soc_videooverlaysoc_record_packetizer_source_last;
assign soc_videooverlaysoc_record_source_source_payload_data = soc_videooverlaysoc_record_packetizer_source_payload_data;
assign soc_videooverlaysoc_record_source_source_payload_error = soc_videooverlaysoc_record_packetizer_source_payload_error;
assign soc_videooverlaysoc_record_source_source_param_addr_size = soc_videooverlaysoc_record_packetizer_source_param_addr_size;
assign soc_videooverlaysoc_record_source_source_param_nr = soc_videooverlaysoc_record_packetizer_source_param_nr;
assign soc_videooverlaysoc_record_source_source_param_pf = soc_videooverlaysoc_record_packetizer_source_param_pf;
assign soc_videooverlaysoc_record_source_source_param_port_size = soc_videooverlaysoc_record_packetizer_source_param_port_size;
assign soc_videooverlaysoc_record_source_source_param_pr = soc_videooverlaysoc_record_packetizer_source_param_pr;
assign soc_videooverlaysoc_record_source_source_param_src_port = soc_videooverlaysoc_record_packetizer_source_param_src_port;
assign soc_videooverlaysoc_record_source_source_param_dst_port = soc_videooverlaysoc_record_packetizer_source_param_dst_port;
always @(*) begin
	soc_videooverlaysoc_record_source_source_param_length <= 16'd0;
	soc_videooverlaysoc_record_source_source_param_length <= soc_videooverlaysoc_record_packetizer_source_param_length;
	soc_videooverlaysoc_record_source_source_param_length <= ((((3'd4 + ((soc_videooverlaysoc_record_sender_source_source_param_wcount != 1'd0) * 3'd4)) + (soc_videooverlaysoc_record_sender_source_source_param_wcount * 3'd4)) + ((soc_videooverlaysoc_record_sender_source_source_param_rcount != 1'd0) * 3'd4)) + (soc_videooverlaysoc_record_sender_source_source_param_rcount * 3'd4));
end
always @(*) begin
	soc_videooverlaysoc_record_source_source_param_ip_address <= 32'd0;
	soc_videooverlaysoc_record_source_source_param_ip_address <= soc_videooverlaysoc_record_packetizer_source_param_ip_address;
	soc_videooverlaysoc_record_source_source_param_ip_address <= soc_videooverlaysoc_record_last_ip_address;
end
always @(*) begin
	soc_videooverlaysoc_record_packetizer_sink_payload_data <= 32'd0;
	soc_videooverlaysoc_record_packetizer_sink_payload_data <= soc_videooverlaysoc_record_sender_source_source_payload_data;
	soc_videooverlaysoc_record_packetizer_sink_payload_data <= {soc_videooverlaysoc_record_sender_source_source_payload_data[7:0], soc_videooverlaysoc_record_sender_source_source_payload_data[15:8], soc_videooverlaysoc_record_sender_source_source_payload_data[23:16], soc_videooverlaysoc_record_sender_source_source_payload_data[31:24]};
end
assign soc_videooverlaysoc_record_depacketizer_header = soc_videooverlaysoc_record_depacketizer_header_reg;
assign soc_videooverlaysoc_record_depacketizer_source_payload_error = soc_videooverlaysoc_record_depacketizer_sink_payload_error;
assign soc_videooverlaysoc_record_depacketizer_source_last = (soc_videooverlaysoc_record_depacketizer_sink_last | soc_videooverlaysoc_record_depacketizer_no_payload);
assign soc_videooverlaysoc_record_depacketizer_source_payload_data = soc_videooverlaysoc_record_depacketizer_sink_payload_data;
assign soc_videooverlaysoc_record_depacketizer_source_param_bca = {vns_slice_proxy84};
assign soc_videooverlaysoc_record_depacketizer_source_param_byte_enable = {vns_slice_proxy85[7:0]};
assign soc_videooverlaysoc_record_depacketizer_source_param_cyc = {vns_slice_proxy86};
assign soc_videooverlaysoc_record_depacketizer_source_param_rca = {vns_slice_proxy87};
assign soc_videooverlaysoc_record_depacketizer_source_param_rcount = {vns_slice_proxy88[7:0]};
assign soc_videooverlaysoc_record_depacketizer_source_param_rff = {vns_slice_proxy89};
assign soc_videooverlaysoc_record_depacketizer_source_param_wca = {vns_slice_proxy90};
assign soc_videooverlaysoc_record_depacketizer_source_param_wcount = {vns_slice_proxy91[7:0]};
assign soc_videooverlaysoc_record_depacketizer_source_param_wff = {vns_slice_proxy92};
always @(*) begin
	soc_videooverlaysoc_record_depacketizer_source_valid <= 1'd0;
	soc_videooverlaysoc_record_depacketizer_shift <= 1'd0;
	vns_liteethetherbonerecorddepacketizer_next_state <= 1'd0;
	soc_videooverlaysoc_record_depacketizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_record_depacketizer_counter_reset <= 1'd0;
	vns_liteethetherbonerecorddepacketizer_next_state <= vns_liteethetherbonerecorddepacketizer_state;
	case (vns_liteethetherbonerecorddepacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_record_depacketizer_sink_ready <= soc_videooverlaysoc_record_depacketizer_source_ready;
			soc_videooverlaysoc_record_depacketizer_source_valid <= (soc_videooverlaysoc_record_depacketizer_sink_valid | soc_videooverlaysoc_record_depacketizer_no_payload);
			if (((soc_videooverlaysoc_record_depacketizer_source_valid & soc_videooverlaysoc_record_depacketizer_source_ready) & soc_videooverlaysoc_record_depacketizer_source_last)) begin
				vns_liteethetherbonerecorddepacketizer_next_state <= 1'd0;
			end
		end
		default: begin
			soc_videooverlaysoc_record_depacketizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_record_depacketizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_record_depacketizer_sink_valid) begin
				soc_videooverlaysoc_record_depacketizer_shift <= 1'd1;
				vns_liteethetherbonerecorddepacketizer_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videooverlaysoc_record_depacketizer_is_el = ((~(vns_liteethetherbonerecorddepacketizer_state == 1'd1)) & (vns_liteethetherbonerecorddepacketizer_next_state == 1'd1));
assign soc_videooverlaysoc_record_receiver_fifo_sink_valid = soc_videooverlaysoc_record_receiver_sink_sink_valid;
assign soc_videooverlaysoc_record_receiver_sink_sink_ready = soc_videooverlaysoc_record_receiver_fifo_sink_ready;
assign soc_videooverlaysoc_record_receiver_fifo_sink_first = soc_videooverlaysoc_record_receiver_sink_sink_first;
assign soc_videooverlaysoc_record_receiver_fifo_sink_last = soc_videooverlaysoc_record_receiver_sink_sink_last;
assign soc_videooverlaysoc_record_receiver_fifo_sink_payload_data = soc_videooverlaysoc_record_receiver_sink_sink_payload_data;
assign soc_videooverlaysoc_record_receiver_fifo_sink_payload_error = soc_videooverlaysoc_record_receiver_sink_sink_payload_error;
assign soc_videooverlaysoc_record_receiver_fifo_sink_param_bca = soc_videooverlaysoc_record_receiver_sink_sink_param_bca;
assign soc_videooverlaysoc_record_receiver_fifo_sink_param_byte_enable = soc_videooverlaysoc_record_receiver_sink_sink_param_byte_enable;
assign soc_videooverlaysoc_record_receiver_fifo_sink_param_cyc = soc_videooverlaysoc_record_receiver_sink_sink_param_cyc;
assign soc_videooverlaysoc_record_receiver_fifo_sink_param_rca = soc_videooverlaysoc_record_receiver_sink_sink_param_rca;
assign soc_videooverlaysoc_record_receiver_fifo_sink_param_rcount = soc_videooverlaysoc_record_receiver_sink_sink_param_rcount;
assign soc_videooverlaysoc_record_receiver_fifo_sink_param_rff = soc_videooverlaysoc_record_receiver_sink_sink_param_rff;
assign soc_videooverlaysoc_record_receiver_fifo_sink_param_wca = soc_videooverlaysoc_record_receiver_sink_sink_param_wca;
assign soc_videooverlaysoc_record_receiver_fifo_sink_param_wcount = soc_videooverlaysoc_record_receiver_sink_sink_param_wcount;
assign soc_videooverlaysoc_record_receiver_fifo_sink_param_wff = soc_videooverlaysoc_record_receiver_sink_sink_param_wff;
assign soc_videooverlaysoc_record_receiver_fifo_syncfifo_din = {soc_videooverlaysoc_record_receiver_fifo_fifo_in_last, soc_videooverlaysoc_record_receiver_fifo_fifo_in_first, soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_wff, soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_wcount, soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_wca, soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_rff, soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_rcount, soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_rca, soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_cyc, soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_byte_enable, soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_bca, soc_videooverlaysoc_record_receiver_fifo_fifo_in_payload_error, soc_videooverlaysoc_record_receiver_fifo_fifo_in_payload_data};
assign {soc_videooverlaysoc_record_receiver_fifo_fifo_out_last, soc_videooverlaysoc_record_receiver_fifo_fifo_out_first, soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_wff, soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_wcount, soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_wca, soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_rff, soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_rcount, soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_rca, soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_cyc, soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_byte_enable, soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_bca, soc_videooverlaysoc_record_receiver_fifo_fifo_out_payload_error, soc_videooverlaysoc_record_receiver_fifo_fifo_out_payload_data} = soc_videooverlaysoc_record_receiver_fifo_syncfifo_dout;
assign soc_videooverlaysoc_record_receiver_fifo_sink_ready = soc_videooverlaysoc_record_receiver_fifo_syncfifo_writable;
assign soc_videooverlaysoc_record_receiver_fifo_syncfifo_we = soc_videooverlaysoc_record_receiver_fifo_sink_valid;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_first = soc_videooverlaysoc_record_receiver_fifo_sink_first;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_last = soc_videooverlaysoc_record_receiver_fifo_sink_last;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_payload_data = soc_videooverlaysoc_record_receiver_fifo_sink_payload_data;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_payload_error = soc_videooverlaysoc_record_receiver_fifo_sink_payload_error;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_bca = soc_videooverlaysoc_record_receiver_fifo_sink_param_bca;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_byte_enable = soc_videooverlaysoc_record_receiver_fifo_sink_param_byte_enable;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_cyc = soc_videooverlaysoc_record_receiver_fifo_sink_param_cyc;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_rca = soc_videooverlaysoc_record_receiver_fifo_sink_param_rca;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_rcount = soc_videooverlaysoc_record_receiver_fifo_sink_param_rcount;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_rff = soc_videooverlaysoc_record_receiver_fifo_sink_param_rff;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_wca = soc_videooverlaysoc_record_receiver_fifo_sink_param_wca;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_wcount = soc_videooverlaysoc_record_receiver_fifo_sink_param_wcount;
assign soc_videooverlaysoc_record_receiver_fifo_fifo_in_param_wff = soc_videooverlaysoc_record_receiver_fifo_sink_param_wff;
assign soc_videooverlaysoc_record_receiver_fifo_source_valid = soc_videooverlaysoc_record_receiver_fifo_readable;
assign soc_videooverlaysoc_record_receiver_fifo_source_first = soc_videooverlaysoc_record_receiver_fifo_fifo_out_first;
assign soc_videooverlaysoc_record_receiver_fifo_source_last = soc_videooverlaysoc_record_receiver_fifo_fifo_out_last;
assign soc_videooverlaysoc_record_receiver_fifo_source_payload_data = soc_videooverlaysoc_record_receiver_fifo_fifo_out_payload_data;
assign soc_videooverlaysoc_record_receiver_fifo_source_payload_error = soc_videooverlaysoc_record_receiver_fifo_fifo_out_payload_error;
assign soc_videooverlaysoc_record_receiver_fifo_source_param_bca = soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_bca;
assign soc_videooverlaysoc_record_receiver_fifo_source_param_byte_enable = soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_byte_enable;
assign soc_videooverlaysoc_record_receiver_fifo_source_param_cyc = soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_cyc;
assign soc_videooverlaysoc_record_receiver_fifo_source_param_rca = soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_rca;
assign soc_videooverlaysoc_record_receiver_fifo_source_param_rcount = soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_rcount;
assign soc_videooverlaysoc_record_receiver_fifo_source_param_rff = soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_rff;
assign soc_videooverlaysoc_record_receiver_fifo_source_param_wca = soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_wca;
assign soc_videooverlaysoc_record_receiver_fifo_source_param_wcount = soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_wcount;
assign soc_videooverlaysoc_record_receiver_fifo_source_param_wff = soc_videooverlaysoc_record_receiver_fifo_fifo_out_param_wff;
assign soc_videooverlaysoc_record_receiver_fifo_re = soc_videooverlaysoc_record_receiver_fifo_source_ready;
assign soc_videooverlaysoc_record_receiver_fifo_syncfifo_re = (soc_videooverlaysoc_record_receiver_fifo_syncfifo_readable & ((~soc_videooverlaysoc_record_receiver_fifo_readable) | soc_videooverlaysoc_record_receiver_fifo_re));
assign soc_videooverlaysoc_record_receiver_fifo_level1 = (soc_videooverlaysoc_record_receiver_fifo_level0 + soc_videooverlaysoc_record_receiver_fifo_readable);
always @(*) begin
	soc_videooverlaysoc_record_receiver_fifo_wrport_adr <= 2'd0;
	if (soc_videooverlaysoc_record_receiver_fifo_replace) begin
		soc_videooverlaysoc_record_receiver_fifo_wrport_adr <= (soc_videooverlaysoc_record_receiver_fifo_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_record_receiver_fifo_wrport_adr <= soc_videooverlaysoc_record_receiver_fifo_produce;
	end
end
assign soc_videooverlaysoc_record_receiver_fifo_wrport_dat_w = soc_videooverlaysoc_record_receiver_fifo_syncfifo_din;
assign soc_videooverlaysoc_record_receiver_fifo_wrport_we = (soc_videooverlaysoc_record_receiver_fifo_syncfifo_we & (soc_videooverlaysoc_record_receiver_fifo_syncfifo_writable | soc_videooverlaysoc_record_receiver_fifo_replace));
assign soc_videooverlaysoc_record_receiver_fifo_do_read = (soc_videooverlaysoc_record_receiver_fifo_syncfifo_readable & soc_videooverlaysoc_record_receiver_fifo_syncfifo_re);
assign soc_videooverlaysoc_record_receiver_fifo_rdport_adr = soc_videooverlaysoc_record_receiver_fifo_consume;
assign soc_videooverlaysoc_record_receiver_fifo_syncfifo_dout = soc_videooverlaysoc_record_receiver_fifo_rdport_dat_r;
assign soc_videooverlaysoc_record_receiver_fifo_rdport_re = soc_videooverlaysoc_record_receiver_fifo_do_read;
assign soc_videooverlaysoc_record_receiver_fifo_syncfifo_writable = (soc_videooverlaysoc_record_receiver_fifo_level0 != 3'd4);
assign soc_videooverlaysoc_record_receiver_fifo_syncfifo_readable = (soc_videooverlaysoc_record_receiver_fifo_level0 != 1'd0);
always @(*) begin
	soc_videooverlaysoc_record_receiver_base_addr_update <= 1'd0;
	soc_videooverlaysoc_record_receiver_source_source_valid <= 1'd0;
	soc_videooverlaysoc_record_receiver_counter_reset <= 1'd0;
	soc_videooverlaysoc_record_receiver_counter_ce <= 1'd0;
	soc_videooverlaysoc_record_receiver_source_source_last <= 1'd0;
	vns_liteethetherbonerecordreceiver_next_state <= 2'd0;
	soc_videooverlaysoc_record_receiver_source_source_payload_addr <= 32'd0;
	soc_videooverlaysoc_record_receiver_source_source_payload_data <= 32'd0;
	soc_videooverlaysoc_record_receiver_source_source_param_we <= 1'd0;
	soc_videooverlaysoc_record_receiver_source_source_param_count <= 8'd0;
	soc_videooverlaysoc_record_receiver_source_source_param_base_addr <= 32'd0;
	soc_videooverlaysoc_record_receiver_source_source_param_be <= 4'd0;
	soc_videooverlaysoc_record_receiver_fifo_source_ready <= 1'd0;
	vns_liteethetherbonerecordreceiver_next_state <= vns_liteethetherbonerecordreceiver_state;
	case (vns_liteethetherbonerecordreceiver_state)
		1'd1: begin
			soc_videooverlaysoc_record_receiver_source_source_valid <= soc_videooverlaysoc_record_receiver_fifo_source_valid;
			soc_videooverlaysoc_record_receiver_source_source_last <= (soc_videooverlaysoc_record_receiver_counter == (soc_videooverlaysoc_record_receiver_fifo_source_param_wcount - 1'd1));
			soc_videooverlaysoc_record_receiver_source_source_param_count <= soc_videooverlaysoc_record_receiver_fifo_source_param_wcount;
			soc_videooverlaysoc_record_receiver_source_source_param_be <= soc_videooverlaysoc_record_receiver_fifo_source_param_byte_enable;
			soc_videooverlaysoc_record_receiver_source_source_payload_addr <= (soc_videooverlaysoc_record_receiver_base_addr[31:2] + soc_videooverlaysoc_record_receiver_counter);
			soc_videooverlaysoc_record_receiver_source_source_param_we <= 1'd1;
			soc_videooverlaysoc_record_receiver_source_source_payload_data <= soc_videooverlaysoc_record_receiver_fifo_source_payload_data;
			soc_videooverlaysoc_record_receiver_fifo_source_ready <= soc_videooverlaysoc_record_receiver_source_source_ready;
			if ((soc_videooverlaysoc_record_receiver_source_source_valid & soc_videooverlaysoc_record_receiver_source_source_ready)) begin
				soc_videooverlaysoc_record_receiver_counter_ce <= 1'd1;
				if (soc_videooverlaysoc_record_receiver_source_source_last) begin
					if (soc_videooverlaysoc_record_receiver_fifo_source_param_rcount) begin
						vns_liteethetherbonerecordreceiver_next_state <= 2'd2;
					end else begin
						vns_liteethetherbonerecordreceiver_next_state <= 1'd0;
					end
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_record_receiver_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_record_receiver_fifo_source_valid) begin
				soc_videooverlaysoc_record_receiver_base_addr_update <= 1'd1;
				vns_liteethetherbonerecordreceiver_next_state <= 2'd3;
			end
		end
		2'd3: begin
			soc_videooverlaysoc_record_receiver_source_source_valid <= soc_videooverlaysoc_record_receiver_fifo_source_valid;
			soc_videooverlaysoc_record_receiver_source_source_last <= (soc_videooverlaysoc_record_receiver_counter == (soc_videooverlaysoc_record_receiver_fifo_source_param_rcount - 1'd1));
			soc_videooverlaysoc_record_receiver_source_source_param_count <= soc_videooverlaysoc_record_receiver_fifo_source_param_rcount;
			soc_videooverlaysoc_record_receiver_source_source_param_base_addr <= soc_videooverlaysoc_record_receiver_base_addr;
			soc_videooverlaysoc_record_receiver_source_source_payload_addr <= soc_videooverlaysoc_record_receiver_fifo_source_payload_data[31:2];
			soc_videooverlaysoc_record_receiver_fifo_source_ready <= soc_videooverlaysoc_record_receiver_source_source_ready;
			if ((soc_videooverlaysoc_record_receiver_source_source_valid & soc_videooverlaysoc_record_receiver_source_source_ready)) begin
				soc_videooverlaysoc_record_receiver_counter_ce <= 1'd1;
				if (soc_videooverlaysoc_record_receiver_source_source_last) begin
					vns_liteethetherbonerecordreceiver_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_record_receiver_fifo_source_ready <= 1'd1;
			soc_videooverlaysoc_record_receiver_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_record_receiver_fifo_source_valid) begin
				soc_videooverlaysoc_record_receiver_base_addr_update <= 1'd1;
				if (soc_videooverlaysoc_record_receiver_fifo_source_param_wcount) begin
					vns_liteethetherbonerecordreceiver_next_state <= 1'd1;
				end else begin
					if (soc_videooverlaysoc_record_receiver_fifo_source_param_rcount) begin
						vns_liteethetherbonerecordreceiver_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_record_sender_fifo_sink_valid = soc_videooverlaysoc_record_sender_sink_sink_valid;
assign soc_videooverlaysoc_record_sender_sink_sink_ready = soc_videooverlaysoc_record_sender_fifo_sink_ready;
assign soc_videooverlaysoc_record_sender_fifo_sink_first = soc_videooverlaysoc_record_sender_sink_sink_first;
assign soc_videooverlaysoc_record_sender_fifo_sink_last = soc_videooverlaysoc_record_sender_sink_sink_last;
assign soc_videooverlaysoc_record_sender_fifo_sink_payload_addr = soc_videooverlaysoc_record_sender_sink_sink_payload_addr;
assign soc_videooverlaysoc_record_sender_fifo_sink_payload_data = soc_videooverlaysoc_record_sender_sink_sink_payload_data;
assign soc_videooverlaysoc_record_sender_fifo_sink_param_we = soc_videooverlaysoc_record_sender_sink_sink_param_we;
assign soc_videooverlaysoc_record_sender_fifo_sink_param_count = soc_videooverlaysoc_record_sender_sink_sink_param_count;
assign soc_videooverlaysoc_record_sender_fifo_sink_param_base_addr = soc_videooverlaysoc_record_sender_sink_sink_param_base_addr;
assign soc_videooverlaysoc_record_sender_fifo_sink_param_be = soc_videooverlaysoc_record_sender_sink_sink_param_be;
assign soc_videooverlaysoc_record_sender_fifo_syncfifo_din = {soc_videooverlaysoc_record_sender_fifo_fifo_in_last, soc_videooverlaysoc_record_sender_fifo_fifo_in_first, soc_videooverlaysoc_record_sender_fifo_fifo_in_param_be, soc_videooverlaysoc_record_sender_fifo_fifo_in_param_base_addr, soc_videooverlaysoc_record_sender_fifo_fifo_in_param_count, soc_videooverlaysoc_record_sender_fifo_fifo_in_param_we, soc_videooverlaysoc_record_sender_fifo_fifo_in_payload_data, soc_videooverlaysoc_record_sender_fifo_fifo_in_payload_addr};
assign {soc_videooverlaysoc_record_sender_fifo_fifo_out_last, soc_videooverlaysoc_record_sender_fifo_fifo_out_first, soc_videooverlaysoc_record_sender_fifo_fifo_out_param_be, soc_videooverlaysoc_record_sender_fifo_fifo_out_param_base_addr, soc_videooverlaysoc_record_sender_fifo_fifo_out_param_count, soc_videooverlaysoc_record_sender_fifo_fifo_out_param_we, soc_videooverlaysoc_record_sender_fifo_fifo_out_payload_data, soc_videooverlaysoc_record_sender_fifo_fifo_out_payload_addr} = soc_videooverlaysoc_record_sender_fifo_syncfifo_dout;
assign soc_videooverlaysoc_record_sender_fifo_sink_ready = soc_videooverlaysoc_record_sender_fifo_syncfifo_writable;
assign soc_videooverlaysoc_record_sender_fifo_syncfifo_we = soc_videooverlaysoc_record_sender_fifo_sink_valid;
assign soc_videooverlaysoc_record_sender_fifo_fifo_in_first = soc_videooverlaysoc_record_sender_fifo_sink_first;
assign soc_videooverlaysoc_record_sender_fifo_fifo_in_last = soc_videooverlaysoc_record_sender_fifo_sink_last;
assign soc_videooverlaysoc_record_sender_fifo_fifo_in_payload_addr = soc_videooverlaysoc_record_sender_fifo_sink_payload_addr;
assign soc_videooverlaysoc_record_sender_fifo_fifo_in_payload_data = soc_videooverlaysoc_record_sender_fifo_sink_payload_data;
assign soc_videooverlaysoc_record_sender_fifo_fifo_in_param_we = soc_videooverlaysoc_record_sender_fifo_sink_param_we;
assign soc_videooverlaysoc_record_sender_fifo_fifo_in_param_count = soc_videooverlaysoc_record_sender_fifo_sink_param_count;
assign soc_videooverlaysoc_record_sender_fifo_fifo_in_param_base_addr = soc_videooverlaysoc_record_sender_fifo_sink_param_base_addr;
assign soc_videooverlaysoc_record_sender_fifo_fifo_in_param_be = soc_videooverlaysoc_record_sender_fifo_sink_param_be;
assign soc_videooverlaysoc_record_sender_fifo_source_valid = soc_videooverlaysoc_record_sender_fifo_readable;
assign soc_videooverlaysoc_record_sender_fifo_source_first = soc_videooverlaysoc_record_sender_fifo_fifo_out_first;
assign soc_videooverlaysoc_record_sender_fifo_source_last = soc_videooverlaysoc_record_sender_fifo_fifo_out_last;
assign soc_videooverlaysoc_record_sender_fifo_source_payload_addr = soc_videooverlaysoc_record_sender_fifo_fifo_out_payload_addr;
assign soc_videooverlaysoc_record_sender_fifo_source_payload_data = soc_videooverlaysoc_record_sender_fifo_fifo_out_payload_data;
assign soc_videooverlaysoc_record_sender_fifo_source_param_we = soc_videooverlaysoc_record_sender_fifo_fifo_out_param_we;
assign soc_videooverlaysoc_record_sender_fifo_source_param_count = soc_videooverlaysoc_record_sender_fifo_fifo_out_param_count;
assign soc_videooverlaysoc_record_sender_fifo_source_param_base_addr = soc_videooverlaysoc_record_sender_fifo_fifo_out_param_base_addr;
assign soc_videooverlaysoc_record_sender_fifo_source_param_be = soc_videooverlaysoc_record_sender_fifo_fifo_out_param_be;
assign soc_videooverlaysoc_record_sender_fifo_re = soc_videooverlaysoc_record_sender_fifo_source_ready;
assign soc_videooverlaysoc_record_sender_fifo_syncfifo_re = (soc_videooverlaysoc_record_sender_fifo_syncfifo_readable & ((~soc_videooverlaysoc_record_sender_fifo_readable) | soc_videooverlaysoc_record_sender_fifo_re));
assign soc_videooverlaysoc_record_sender_fifo_level1 = (soc_videooverlaysoc_record_sender_fifo_level0 + soc_videooverlaysoc_record_sender_fifo_readable);
always @(*) begin
	soc_videooverlaysoc_record_sender_fifo_wrport_adr <= 2'd0;
	if (soc_videooverlaysoc_record_sender_fifo_replace) begin
		soc_videooverlaysoc_record_sender_fifo_wrport_adr <= (soc_videooverlaysoc_record_sender_fifo_produce - 1'd1);
	end else begin
		soc_videooverlaysoc_record_sender_fifo_wrport_adr <= soc_videooverlaysoc_record_sender_fifo_produce;
	end
end
assign soc_videooverlaysoc_record_sender_fifo_wrport_dat_w = soc_videooverlaysoc_record_sender_fifo_syncfifo_din;
assign soc_videooverlaysoc_record_sender_fifo_wrport_we = (soc_videooverlaysoc_record_sender_fifo_syncfifo_we & (soc_videooverlaysoc_record_sender_fifo_syncfifo_writable | soc_videooverlaysoc_record_sender_fifo_replace));
assign soc_videooverlaysoc_record_sender_fifo_do_read = (soc_videooverlaysoc_record_sender_fifo_syncfifo_readable & soc_videooverlaysoc_record_sender_fifo_syncfifo_re);
assign soc_videooverlaysoc_record_sender_fifo_rdport_adr = soc_videooverlaysoc_record_sender_fifo_consume;
assign soc_videooverlaysoc_record_sender_fifo_syncfifo_dout = soc_videooverlaysoc_record_sender_fifo_rdport_dat_r;
assign soc_videooverlaysoc_record_sender_fifo_rdport_re = soc_videooverlaysoc_record_sender_fifo_do_read;
assign soc_videooverlaysoc_record_sender_fifo_syncfifo_writable = (soc_videooverlaysoc_record_sender_fifo_level0 != 3'd4);
assign soc_videooverlaysoc_record_sender_fifo_syncfifo_readable = (soc_videooverlaysoc_record_sender_fifo_level0 != 1'd0);
always @(*) begin
	soc_videooverlaysoc_record_sender_fifo_source_ready <= 1'd0;
	soc_videooverlaysoc_record_sender_source_source_last <= 1'd0;
	vns_liteethetherbonerecordsender_next_state <= 2'd0;
	soc_videooverlaysoc_record_sender_data_sel <= 1'd0;
	soc_videooverlaysoc_record_sender_source_source_valid <= 1'd0;
	vns_liteethetherbonerecordsender_next_state <= vns_liteethetherbonerecordsender_state;
	case (vns_liteethetherbonerecordsender_state)
		1'd1: begin
			soc_videooverlaysoc_record_sender_source_source_valid <= 1'd1;
			soc_videooverlaysoc_record_sender_source_source_last <= 1'd0;
			if (soc_videooverlaysoc_record_sender_source_source_ready) begin
				soc_videooverlaysoc_record_sender_data_sel <= 1'd1;
				vns_liteethetherbonerecordsender_next_state <= 2'd2;
			end
		end
		2'd2: begin
			soc_videooverlaysoc_record_sender_source_source_valid <= 1'd1;
			soc_videooverlaysoc_record_sender_source_source_last <= soc_videooverlaysoc_record_sender_fifo_source_last;
			soc_videooverlaysoc_record_sender_data_sel <= 1'd1;
			if ((soc_videooverlaysoc_record_sender_source_source_valid & soc_videooverlaysoc_record_sender_source_source_ready)) begin
				soc_videooverlaysoc_record_sender_fifo_source_ready <= 1'd1;
				if (soc_videooverlaysoc_record_sender_source_source_last) begin
					vns_liteethetherbonerecordsender_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_record_sender_fifo_source_ready <= 1'd1;
			if (soc_videooverlaysoc_record_sender_fifo_source_valid) begin
				soc_videooverlaysoc_record_sender_fifo_source_ready <= 1'd0;
				vns_liteethetherbonerecordsender_next_state <= 1'd1;
			end
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_record_packetizer_header <= 32'd0;
	soc_videooverlaysoc_record_packetizer_header[0] <= {soc_videooverlaysoc_record_packetizer_sink_param_bca};
	soc_videooverlaysoc_record_packetizer_header[15:8] <= {soc_videooverlaysoc_record_packetizer_sink_param_byte_enable[7:0]};
	soc_videooverlaysoc_record_packetizer_header[4] <= {soc_videooverlaysoc_record_packetizer_sink_param_cyc};
	soc_videooverlaysoc_record_packetizer_header[1] <= {soc_videooverlaysoc_record_packetizer_sink_param_rca};
	soc_videooverlaysoc_record_packetizer_header[31:24] <= {soc_videooverlaysoc_record_packetizer_sink_param_rcount[7:0]};
	soc_videooverlaysoc_record_packetizer_header[2] <= {soc_videooverlaysoc_record_packetizer_sink_param_rff};
	soc_videooverlaysoc_record_packetizer_header[5] <= {soc_videooverlaysoc_record_packetizer_sink_param_wca};
	soc_videooverlaysoc_record_packetizer_header[23:16] <= {soc_videooverlaysoc_record_packetizer_sink_param_wcount[7:0]};
	soc_videooverlaysoc_record_packetizer_header[6] <= {soc_videooverlaysoc_record_packetizer_sink_param_wff};
end
assign soc_videooverlaysoc_record_packetizer_source_payload_error = soc_videooverlaysoc_record_packetizer_sink_payload_error;
always @(*) begin
	vns_liteethetherbonerecordpacketizer_next_state <= 1'd0;
	soc_videooverlaysoc_record_packetizer_source_valid <= 1'd0;
	soc_videooverlaysoc_record_packetizer_counter_reset <= 1'd0;
	soc_videooverlaysoc_record_packetizer_load <= 1'd0;
	soc_videooverlaysoc_record_packetizer_sink_ready <= 1'd0;
	soc_videooverlaysoc_record_packetizer_source_last <= 1'd0;
	soc_videooverlaysoc_record_packetizer_source_payload_data <= 32'd0;
	vns_liteethetherbonerecordpacketizer_next_state <= vns_liteethetherbonerecordpacketizer_state;
	case (vns_liteethetherbonerecordpacketizer_state)
		1'd1: begin
			soc_videooverlaysoc_record_packetizer_source_valid <= soc_videooverlaysoc_record_packetizer_sink_valid;
			soc_videooverlaysoc_record_packetizer_source_last <= soc_videooverlaysoc_record_packetizer_sink_last;
			soc_videooverlaysoc_record_packetizer_source_payload_data <= soc_videooverlaysoc_record_packetizer_sink_payload_data;
			if ((soc_videooverlaysoc_record_packetizer_source_valid & soc_videooverlaysoc_record_packetizer_source_ready)) begin
				soc_videooverlaysoc_record_packetizer_sink_ready <= 1'd1;
				if (soc_videooverlaysoc_record_packetizer_source_last) begin
					vns_liteethetherbonerecordpacketizer_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_record_packetizer_sink_ready <= 1'd1;
			soc_videooverlaysoc_record_packetizer_counter_reset <= 1'd1;
			if (soc_videooverlaysoc_record_packetizer_sink_valid) begin
				soc_videooverlaysoc_record_packetizer_sink_ready <= 1'd0;
				soc_videooverlaysoc_record_packetizer_source_valid <= 1'd1;
				soc_videooverlaysoc_record_packetizer_source_last <= 1'd0;
				soc_videooverlaysoc_record_packetizer_source_payload_data <= soc_videooverlaysoc_record_packetizer_header[31:0];
				if ((soc_videooverlaysoc_record_packetizer_source_valid & soc_videooverlaysoc_record_packetizer_source_ready)) begin
					soc_videooverlaysoc_record_packetizer_load <= 1'd1;
					vns_liteethetherbonerecordpacketizer_next_state <= 1'd1;
				end
			end
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_dispatcher_sel1 <= 1'd0;
	if (soc_videooverlaysoc_dispatcher_first) begin
		soc_videooverlaysoc_dispatcher_sel1 <= soc_videooverlaysoc_dispatcher_sel0;
	end else begin
		soc_videooverlaysoc_dispatcher_sel1 <= soc_videooverlaysoc_dispatcher_sel_ongoing;
	end
end
always @(*) begin
	soc_videooverlaysoc_packet_source_source_ready <= 1'd0;
	soc_videooverlaysoc_probe_sink_valid <= 1'd0;
	soc_videooverlaysoc_record_sink_sink_valid <= 1'd0;
	soc_videooverlaysoc_probe_sink_first <= 1'd0;
	soc_videooverlaysoc_record_sink_sink_first <= 1'd0;
	soc_videooverlaysoc_probe_sink_last <= 1'd0;
	soc_videooverlaysoc_record_sink_sink_last <= 1'd0;
	soc_videooverlaysoc_probe_sink_payload_data <= 32'd0;
	soc_videooverlaysoc_record_sink_sink_payload_data <= 32'd0;
	soc_videooverlaysoc_probe_sink_payload_error <= 4'd0;
	soc_videooverlaysoc_record_sink_sink_payload_error <= 4'd0;
	soc_videooverlaysoc_probe_sink_param_addr_size <= 4'd0;
	soc_videooverlaysoc_record_sink_sink_param_addr_size <= 4'd0;
	soc_videooverlaysoc_probe_sink_param_nr <= 1'd0;
	soc_videooverlaysoc_record_sink_sink_param_nr <= 1'd0;
	soc_videooverlaysoc_probe_sink_param_pf <= 1'd0;
	soc_videooverlaysoc_record_sink_sink_param_pf <= 1'd0;
	soc_videooverlaysoc_probe_sink_param_port_size <= 4'd0;
	soc_videooverlaysoc_record_sink_sink_param_port_size <= 4'd0;
	soc_videooverlaysoc_probe_sink_param_pr <= 1'd0;
	soc_videooverlaysoc_record_sink_sink_param_pr <= 1'd0;
	soc_videooverlaysoc_probe_sink_param_src_port <= 16'd0;
	soc_videooverlaysoc_record_sink_sink_param_src_port <= 16'd0;
	soc_videooverlaysoc_probe_sink_param_dst_port <= 16'd0;
	soc_videooverlaysoc_record_sink_sink_param_dst_port <= 16'd0;
	soc_videooverlaysoc_probe_sink_param_ip_address <= 32'd0;
	soc_videooverlaysoc_record_sink_sink_param_ip_address <= 32'd0;
	soc_videooverlaysoc_probe_sink_param_length <= 16'd0;
	soc_videooverlaysoc_record_sink_sink_param_length <= 16'd0;
	case (soc_videooverlaysoc_dispatcher_sel1)
		1'd0: begin
			soc_videooverlaysoc_probe_sink_valid <= soc_videooverlaysoc_packet_source_source_valid;
			soc_videooverlaysoc_packet_source_source_ready <= soc_videooverlaysoc_probe_sink_ready;
			soc_videooverlaysoc_probe_sink_first <= soc_videooverlaysoc_packet_source_source_first;
			soc_videooverlaysoc_probe_sink_last <= soc_videooverlaysoc_packet_source_source_last;
			soc_videooverlaysoc_probe_sink_payload_data <= soc_videooverlaysoc_packet_source_source_payload_data;
			soc_videooverlaysoc_probe_sink_payload_error <= soc_videooverlaysoc_packet_source_source_payload_error;
			soc_videooverlaysoc_probe_sink_param_addr_size <= soc_videooverlaysoc_packet_source_source_param_addr_size;
			soc_videooverlaysoc_probe_sink_param_nr <= soc_videooverlaysoc_packet_source_source_param_nr;
			soc_videooverlaysoc_probe_sink_param_pf <= soc_videooverlaysoc_packet_source_source_param_pf;
			soc_videooverlaysoc_probe_sink_param_port_size <= soc_videooverlaysoc_packet_source_source_param_port_size;
			soc_videooverlaysoc_probe_sink_param_pr <= soc_videooverlaysoc_packet_source_source_param_pr;
			soc_videooverlaysoc_probe_sink_param_src_port <= soc_videooverlaysoc_packet_source_source_param_src_port;
			soc_videooverlaysoc_probe_sink_param_dst_port <= soc_videooverlaysoc_packet_source_source_param_dst_port;
			soc_videooverlaysoc_probe_sink_param_ip_address <= soc_videooverlaysoc_packet_source_source_param_ip_address;
			soc_videooverlaysoc_probe_sink_param_length <= soc_videooverlaysoc_packet_source_source_param_length;
		end
		1'd1: begin
			soc_videooverlaysoc_record_sink_sink_valid <= soc_videooverlaysoc_packet_source_source_valid;
			soc_videooverlaysoc_packet_source_source_ready <= soc_videooverlaysoc_record_sink_sink_ready;
			soc_videooverlaysoc_record_sink_sink_first <= soc_videooverlaysoc_packet_source_source_first;
			soc_videooverlaysoc_record_sink_sink_last <= soc_videooverlaysoc_packet_source_source_last;
			soc_videooverlaysoc_record_sink_sink_payload_data <= soc_videooverlaysoc_packet_source_source_payload_data;
			soc_videooverlaysoc_record_sink_sink_payload_error <= soc_videooverlaysoc_packet_source_source_payload_error;
			soc_videooverlaysoc_record_sink_sink_param_addr_size <= soc_videooverlaysoc_packet_source_source_param_addr_size;
			soc_videooverlaysoc_record_sink_sink_param_nr <= soc_videooverlaysoc_packet_source_source_param_nr;
			soc_videooverlaysoc_record_sink_sink_param_pf <= soc_videooverlaysoc_packet_source_source_param_pf;
			soc_videooverlaysoc_record_sink_sink_param_port_size <= soc_videooverlaysoc_packet_source_source_param_port_size;
			soc_videooverlaysoc_record_sink_sink_param_pr <= soc_videooverlaysoc_packet_source_source_param_pr;
			soc_videooverlaysoc_record_sink_sink_param_src_port <= soc_videooverlaysoc_packet_source_source_param_src_port;
			soc_videooverlaysoc_record_sink_sink_param_dst_port <= soc_videooverlaysoc_packet_source_source_param_dst_port;
			soc_videooverlaysoc_record_sink_sink_param_ip_address <= soc_videooverlaysoc_packet_source_source_param_ip_address;
			soc_videooverlaysoc_record_sink_sink_param_length <= soc_videooverlaysoc_packet_source_source_param_length;
		end
		default: begin
			soc_videooverlaysoc_packet_source_source_ready <= 1'd1;
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_dispatcher_last <= 1'd0;
	if (soc_videooverlaysoc_packet_source_source_valid) begin
		soc_videooverlaysoc_dispatcher_last <= (soc_videooverlaysoc_packet_source_source_last & soc_videooverlaysoc_packet_source_source_ready);
	end
end
assign soc_videooverlaysoc_dispatcher_ongoing0 = ((soc_videooverlaysoc_packet_source_source_valid | soc_videooverlaysoc_dispatcher_ongoing1) & (~soc_videooverlaysoc_dispatcher_last));
always @(*) begin
	soc_videooverlaysoc_request <= 2'd0;
	soc_videooverlaysoc_request[0] <= soc_videooverlaysoc_status0_ongoing0;
	soc_videooverlaysoc_request[1] <= soc_videooverlaysoc_status1_ongoing0;
end
always @(*) begin
	soc_videooverlaysoc_packet_sink_valid <= 1'd0;
	soc_videooverlaysoc_packet_sink_first <= 1'd0;
	soc_videooverlaysoc_packet_sink_last <= 1'd0;
	soc_videooverlaysoc_packet_sink_payload_data <= 32'd0;
	soc_videooverlaysoc_packet_sink_payload_error <= 4'd0;
	soc_videooverlaysoc_packet_sink_param_addr_size <= 4'd0;
	soc_videooverlaysoc_packet_sink_param_nr <= 1'd0;
	soc_videooverlaysoc_packet_sink_param_pf <= 1'd0;
	soc_videooverlaysoc_packet_sink_param_port_size <= 4'd0;
	soc_videooverlaysoc_packet_sink_param_pr <= 1'd0;
	soc_videooverlaysoc_packet_sink_param_src_port <= 16'd0;
	soc_videooverlaysoc_packet_sink_param_dst_port <= 16'd0;
	soc_videooverlaysoc_packet_sink_param_ip_address <= 32'd0;
	soc_videooverlaysoc_packet_sink_param_length <= 16'd0;
	soc_videooverlaysoc_probe_source_ready <= 1'd0;
	soc_videooverlaysoc_record_source_source_ready <= 1'd0;
	case (soc_videooverlaysoc_grant)
		1'd0: begin
			soc_videooverlaysoc_packet_sink_valid <= soc_videooverlaysoc_probe_source_valid;
			soc_videooverlaysoc_probe_source_ready <= soc_videooverlaysoc_packet_sink_ready;
			soc_videooverlaysoc_packet_sink_first <= soc_videooverlaysoc_probe_source_first;
			soc_videooverlaysoc_packet_sink_last <= soc_videooverlaysoc_probe_source_last;
			soc_videooverlaysoc_packet_sink_payload_data <= soc_videooverlaysoc_probe_source_payload_data;
			soc_videooverlaysoc_packet_sink_payload_error <= soc_videooverlaysoc_probe_source_payload_error;
			soc_videooverlaysoc_packet_sink_param_addr_size <= soc_videooverlaysoc_probe_source_param_addr_size;
			soc_videooverlaysoc_packet_sink_param_nr <= soc_videooverlaysoc_probe_source_param_nr;
			soc_videooverlaysoc_packet_sink_param_pf <= soc_videooverlaysoc_probe_source_param_pf;
			soc_videooverlaysoc_packet_sink_param_port_size <= soc_videooverlaysoc_probe_source_param_port_size;
			soc_videooverlaysoc_packet_sink_param_pr <= soc_videooverlaysoc_probe_source_param_pr;
			soc_videooverlaysoc_packet_sink_param_src_port <= soc_videooverlaysoc_probe_source_param_src_port;
			soc_videooverlaysoc_packet_sink_param_dst_port <= soc_videooverlaysoc_probe_source_param_dst_port;
			soc_videooverlaysoc_packet_sink_param_ip_address <= soc_videooverlaysoc_probe_source_param_ip_address;
			soc_videooverlaysoc_packet_sink_param_length <= soc_videooverlaysoc_probe_source_param_length;
		end
		1'd1: begin
			soc_videooverlaysoc_packet_sink_valid <= soc_videooverlaysoc_record_source_source_valid;
			soc_videooverlaysoc_record_source_source_ready <= soc_videooverlaysoc_packet_sink_ready;
			soc_videooverlaysoc_packet_sink_first <= soc_videooverlaysoc_record_source_source_first;
			soc_videooverlaysoc_packet_sink_last <= soc_videooverlaysoc_record_source_source_last;
			soc_videooverlaysoc_packet_sink_payload_data <= soc_videooverlaysoc_record_source_source_payload_data;
			soc_videooverlaysoc_packet_sink_payload_error <= soc_videooverlaysoc_record_source_source_payload_error;
			soc_videooverlaysoc_packet_sink_param_addr_size <= soc_videooverlaysoc_record_source_source_param_addr_size;
			soc_videooverlaysoc_packet_sink_param_nr <= soc_videooverlaysoc_record_source_source_param_nr;
			soc_videooverlaysoc_packet_sink_param_pf <= soc_videooverlaysoc_record_source_source_param_pf;
			soc_videooverlaysoc_packet_sink_param_port_size <= soc_videooverlaysoc_record_source_source_param_port_size;
			soc_videooverlaysoc_packet_sink_param_pr <= soc_videooverlaysoc_record_source_source_param_pr;
			soc_videooverlaysoc_packet_sink_param_src_port <= soc_videooverlaysoc_record_source_source_param_src_port;
			soc_videooverlaysoc_packet_sink_param_dst_port <= soc_videooverlaysoc_record_source_source_param_dst_port;
			soc_videooverlaysoc_packet_sink_param_ip_address <= soc_videooverlaysoc_record_source_source_param_ip_address;
			soc_videooverlaysoc_packet_sink_param_length <= soc_videooverlaysoc_record_source_source_param_length;
		end
	endcase
end
always @(*) begin
	soc_videooverlaysoc_status0_last <= 1'd0;
	if (soc_videooverlaysoc_probe_source_valid) begin
		soc_videooverlaysoc_status0_last <= (soc_videooverlaysoc_probe_source_last & soc_videooverlaysoc_probe_source_ready);
	end
end
assign soc_videooverlaysoc_status0_ongoing0 = ((soc_videooverlaysoc_probe_source_valid | soc_videooverlaysoc_status0_ongoing1) & (~soc_videooverlaysoc_status0_last));
always @(*) begin
	soc_videooverlaysoc_status1_last <= 1'd0;
	if (soc_videooverlaysoc_record_source_source_valid) begin
		soc_videooverlaysoc_status1_last <= (soc_videooverlaysoc_record_source_source_last & soc_videooverlaysoc_record_source_source_ready);
	end
end
assign soc_videooverlaysoc_status1_ongoing0 = ((soc_videooverlaysoc_record_source_source_valid | soc_videooverlaysoc_status1_ongoing1) & (~soc_videooverlaysoc_status1_last));
always @(*) begin
	soc_videooverlaysoc_wishbone_sink_ready <= 1'd0;
	soc_videooverlaysoc_wishbone_bus_adr <= 30'd0;
	soc_videooverlaysoc_wishbone_bus_dat_w <= 32'd0;
	soc_videooverlaysoc_wishbone_bus_sel <= 4'd0;
	soc_videooverlaysoc_wishbone_bus_cyc <= 1'd0;
	soc_videooverlaysoc_wishbone_bus_stb <= 1'd0;
	soc_videooverlaysoc_wishbone_source_valid <= 1'd0;
	soc_videooverlaysoc_wishbone_bus_we <= 1'd0;
	soc_videooverlaysoc_wishbone_source_last <= 1'd0;
	soc_videooverlaysoc_wishbone_data_update <= 1'd0;
	vns_liteethetherbonewishbonemaster_next_state <= 2'd0;
	vns_liteethetherbonewishbonemaster_next_state <= vns_liteethetherbonewishbonemaster_state;
	case (vns_liteethetherbonewishbonemaster_state)
		1'd1: begin
			soc_videooverlaysoc_wishbone_bus_adr <= soc_videooverlaysoc_wishbone_sink_payload_addr;
			soc_videooverlaysoc_wishbone_bus_dat_w <= soc_videooverlaysoc_wishbone_sink_payload_data;
			soc_videooverlaysoc_wishbone_bus_sel <= soc_videooverlaysoc_wishbone_sink_param_be;
			soc_videooverlaysoc_wishbone_bus_stb <= soc_videooverlaysoc_wishbone_sink_valid;
			soc_videooverlaysoc_wishbone_bus_we <= 1'd1;
			soc_videooverlaysoc_wishbone_bus_cyc <= 1'd1;
			if ((soc_videooverlaysoc_wishbone_bus_stb & soc_videooverlaysoc_wishbone_bus_ack)) begin
				soc_videooverlaysoc_wishbone_sink_ready <= 1'd1;
				if (soc_videooverlaysoc_wishbone_sink_last) begin
					vns_liteethetherbonewishbonemaster_next_state <= 1'd0;
				end
			end
		end
		2'd2: begin
			soc_videooverlaysoc_wishbone_bus_adr <= soc_videooverlaysoc_wishbone_sink_payload_addr;
			soc_videooverlaysoc_wishbone_bus_sel <= soc_videooverlaysoc_wishbone_sink_param_be;
			soc_videooverlaysoc_wishbone_bus_stb <= soc_videooverlaysoc_wishbone_sink_valid;
			soc_videooverlaysoc_wishbone_bus_cyc <= 1'd1;
			if ((soc_videooverlaysoc_wishbone_bus_stb & soc_videooverlaysoc_wishbone_bus_ack)) begin
				soc_videooverlaysoc_wishbone_data_update <= 1'd1;
				vns_liteethetherbonewishbonemaster_next_state <= 2'd3;
			end
		end
		2'd3: begin
			soc_videooverlaysoc_wishbone_source_valid <= soc_videooverlaysoc_wishbone_sink_valid;
			soc_videooverlaysoc_wishbone_source_last <= soc_videooverlaysoc_wishbone_sink_last;
			if ((soc_videooverlaysoc_wishbone_source_valid & soc_videooverlaysoc_wishbone_source_ready)) begin
				soc_videooverlaysoc_wishbone_sink_ready <= 1'd1;
				if (soc_videooverlaysoc_wishbone_source_last) begin
					vns_liteethetherbonewishbonemaster_next_state <= 1'd0;
				end else begin
					vns_liteethetherbonewishbonemaster_next_state <= 2'd2;
				end
			end
		end
		default: begin
			soc_videooverlaysoc_wishbone_sink_ready <= 1'd1;
			if (soc_videooverlaysoc_wishbone_sink_valid) begin
				soc_videooverlaysoc_wishbone_sink_ready <= 1'd0;
				if (soc_videooverlaysoc_wishbone_sink_param_we) begin
					vns_liteethetherbonewishbonemaster_next_state <= 1'd1;
				end else begin
					vns_liteethetherbonewishbonemaster_next_state <= 2'd2;
				end
			end
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr = vns_comb_rhs_array_muxed38;
assign soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_w = vns_comb_rhs_array_muxed39;
assign soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_sel = vns_comb_rhs_array_muxed40;
assign soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_cyc = vns_comb_rhs_array_muxed41;
assign soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_stb = vns_comb_rhs_array_muxed42;
assign soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_we = vns_comb_rhs_array_muxed43;
assign soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_cti = vns_comb_rhs_array_muxed44;
assign soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_bte = vns_comb_rhs_array_muxed45;
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_dat_r = soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_ack = (soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_ack & (vns_wb_sdram_con_grant == 1'd0));
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_err = (soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_err & (vns_wb_sdram_con_grant == 1'd0));
assign vns_wb_sdram_con_request = {soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_cyc};
assign vns_wb_sdram_con_grant = 1'd0;
assign vns_videooverlaysoc_shared_adr = vns_comb_rhs_array_muxed46;
assign vns_videooverlaysoc_shared_dat_w = vns_comb_rhs_array_muxed47;
assign vns_videooverlaysoc_shared_sel = vns_comb_rhs_array_muxed48;
assign vns_videooverlaysoc_shared_cyc = vns_comb_rhs_array_muxed49;
assign vns_videooverlaysoc_shared_stb = vns_comb_rhs_array_muxed50;
assign vns_videooverlaysoc_shared_we = vns_comb_rhs_array_muxed51;
assign vns_videooverlaysoc_shared_cti = vns_comb_rhs_array_muxed52;
assign vns_videooverlaysoc_shared_bte = vns_comb_rhs_array_muxed53;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_dat_r = vns_videooverlaysoc_shared_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_dat_r = vns_videooverlaysoc_shared_dat_r;
assign soc_videooverlaysoc_wishbone_bus_dat_r = vns_videooverlaysoc_shared_dat_r;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_ack = (vns_videooverlaysoc_shared_ack & (vns_videooverlaysoc_grant == 1'd0));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_ack = (vns_videooverlaysoc_shared_ack & (vns_videooverlaysoc_grant == 1'd1));
assign soc_videooverlaysoc_wishbone_bus_ack = (vns_videooverlaysoc_shared_ack & (vns_videooverlaysoc_grant == 2'd2));
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_err <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_err <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_err;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_err <= (vns_videooverlaysoc_shared_err & (vns_videooverlaysoc_grant == 1'd0));
end
always @(*) begin
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_err <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_err <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_d_err;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_err <= (vns_videooverlaysoc_shared_err & (vns_videooverlaysoc_grant == 1'd1));
end
assign soc_videooverlaysoc_wishbone_bus_err = (vns_videooverlaysoc_shared_err & (vns_videooverlaysoc_grant == 2'd2));
assign vns_videooverlaysoc_request = {soc_videooverlaysoc_wishbone_bus_cyc, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_cyc, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_cyc};
always @(*) begin
	vns_videooverlaysoc_slave_sel <= 5'd0;
	vns_videooverlaysoc_slave_sel[0] <= (vns_videooverlaysoc_shared_adr[28:26] == 1'd0);
	vns_videooverlaysoc_slave_sel[1] <= (vns_videooverlaysoc_shared_adr[28:26] == 1'd1);
	vns_videooverlaysoc_slave_sel[2] <= (vns_videooverlaysoc_shared_adr[28:26] == 3'd6);
	vns_videooverlaysoc_slave_sel[3] <= (vns_videooverlaysoc_shared_adr[28:26] == 3'd4);
	vns_videooverlaysoc_slave_sel[4] <= (vns_videooverlaysoc_shared_adr[28:26] == 3'd7);
end
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_adr = vns_videooverlaysoc_shared_adr;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_dat_w = vns_videooverlaysoc_shared_dat_w;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_sel = vns_videooverlaysoc_shared_sel;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_stb = vns_videooverlaysoc_shared_stb;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_we = vns_videooverlaysoc_shared_we;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_cti = vns_videooverlaysoc_shared_cti;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_bte = vns_videooverlaysoc_shared_bte;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_adr = vns_videooverlaysoc_shared_adr;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_dat_w = vns_videooverlaysoc_shared_dat_w;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_sel = vns_videooverlaysoc_shared_sel;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_stb = vns_videooverlaysoc_shared_stb;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_we = vns_videooverlaysoc_shared_we;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_cti = vns_videooverlaysoc_shared_cti;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_bte = vns_videooverlaysoc_shared_bte;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_adr = vns_videooverlaysoc_shared_adr;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_dat_w = vns_videooverlaysoc_shared_dat_w;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_sel = vns_videooverlaysoc_shared_sel;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_stb = vns_videooverlaysoc_shared_stb;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_we = vns_videooverlaysoc_shared_we;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_cti = vns_videooverlaysoc_shared_cti;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_bte = vns_videooverlaysoc_shared_bte;
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_adr = vns_videooverlaysoc_shared_adr;
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_dat_w = vns_videooverlaysoc_shared_dat_w;
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_sel = vns_videooverlaysoc_shared_sel;
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_stb = vns_videooverlaysoc_shared_stb;
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_we = vns_videooverlaysoc_shared_we;
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_cti = vns_videooverlaysoc_shared_cti;
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_bte = vns_videooverlaysoc_shared_bte;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_adr = vns_videooverlaysoc_shared_adr;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_dat_w = vns_videooverlaysoc_shared_dat_w;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_sel = vns_videooverlaysoc_shared_sel;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_stb = vns_videooverlaysoc_shared_stb;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_we = vns_videooverlaysoc_shared_we;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_cti = vns_videooverlaysoc_shared_cti;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_bte = vns_videooverlaysoc_shared_bte;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_cyc = (vns_videooverlaysoc_shared_cyc & vns_videooverlaysoc_slave_sel[0]);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_cyc = (vns_videooverlaysoc_shared_cyc & vns_videooverlaysoc_slave_sel[1]);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_cyc = (vns_videooverlaysoc_shared_cyc & vns_videooverlaysoc_slave_sel[2]);
assign soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_cyc = (vns_videooverlaysoc_shared_cyc & vns_videooverlaysoc_slave_sel[3]);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_cyc = (vns_videooverlaysoc_shared_cyc & vns_videooverlaysoc_slave_sel[4]);
assign vns_videooverlaysoc_shared_err = ((((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_err | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_err) | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_err) | soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_err) | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_err);
assign vns_videooverlaysoc_wait = ((vns_videooverlaysoc_shared_stb & vns_videooverlaysoc_shared_cyc) & (~vns_videooverlaysoc_shared_ack));
always @(*) begin
	vns_videooverlaysoc_shared_dat_r <= 32'd0;
	vns_videooverlaysoc_shared_ack <= 1'd0;
	vns_videooverlaysoc_error <= 1'd0;
	vns_videooverlaysoc_shared_ack <= ((((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_ack | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_ack) | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_ack) | soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_ack) | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_ack);
	vns_videooverlaysoc_shared_dat_r <= ((((({32{vns_videooverlaysoc_slave_sel_r[0]}} & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_dat_r) | ({32{vns_videooverlaysoc_slave_sel_r[1]}} & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_dat_r)) | ({32{vns_videooverlaysoc_slave_sel_r[2]}} & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_dat_r)) | ({32{vns_videooverlaysoc_slave_sel_r[3]}} & soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_dat_r)) | ({32{vns_videooverlaysoc_slave_sel_r[4]}} & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_dat_r));
	if (vns_videooverlaysoc_done) begin
		vns_videooverlaysoc_shared_dat_r <= 32'd4294967295;
		vns_videooverlaysoc_shared_ack <= 1'd1;
		vns_videooverlaysoc_error <= 1'd1;
	end
end
assign vns_videooverlaysoc_done = (vns_videooverlaysoc_count == 1'd0);
assign vns_videooverlaysoc_csrbank0_sel = (vns_videooverlaysoc_interface0_bank_bus_adr[13:9] == 1'd0);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_reset_reset_r = vns_videooverlaysoc_interface0_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_reset_reset_re = ((vns_videooverlaysoc_csrbank0_sel & vns_videooverlaysoc_interface0_bank_bus_we) & (vns_videooverlaysoc_interface0_bank_bus_adr[3:0] == 1'd0));
assign vns_videooverlaysoc_csrbank0_scratch3_r = vns_videooverlaysoc_interface0_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank0_scratch3_re = ((vns_videooverlaysoc_csrbank0_sel & vns_videooverlaysoc_interface0_bank_bus_we) & (vns_videooverlaysoc_interface0_bank_bus_adr[3:0] == 1'd1));
assign vns_videooverlaysoc_csrbank0_scratch2_r = vns_videooverlaysoc_interface0_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank0_scratch2_re = ((vns_videooverlaysoc_csrbank0_sel & vns_videooverlaysoc_interface0_bank_bus_we) & (vns_videooverlaysoc_interface0_bank_bus_adr[3:0] == 2'd2));
assign vns_videooverlaysoc_csrbank0_scratch1_r = vns_videooverlaysoc_interface0_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank0_scratch1_re = ((vns_videooverlaysoc_csrbank0_sel & vns_videooverlaysoc_interface0_bank_bus_we) & (vns_videooverlaysoc_interface0_bank_bus_adr[3:0] == 2'd3));
assign vns_videooverlaysoc_csrbank0_scratch0_r = vns_videooverlaysoc_interface0_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank0_scratch0_re = ((vns_videooverlaysoc_csrbank0_sel & vns_videooverlaysoc_interface0_bank_bus_we) & (vns_videooverlaysoc_interface0_bank_bus_adr[3:0] == 3'd4));
assign vns_videooverlaysoc_csrbank0_bus_errors3_r = vns_videooverlaysoc_interface0_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank0_bus_errors3_re = ((vns_videooverlaysoc_csrbank0_sel & vns_videooverlaysoc_interface0_bank_bus_we) & (vns_videooverlaysoc_interface0_bank_bus_adr[3:0] == 3'd5));
assign vns_videooverlaysoc_csrbank0_bus_errors2_r = vns_videooverlaysoc_interface0_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank0_bus_errors2_re = ((vns_videooverlaysoc_csrbank0_sel & vns_videooverlaysoc_interface0_bank_bus_we) & (vns_videooverlaysoc_interface0_bank_bus_adr[3:0] == 3'd6));
assign vns_videooverlaysoc_csrbank0_bus_errors1_r = vns_videooverlaysoc_interface0_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank0_bus_errors1_re = ((vns_videooverlaysoc_csrbank0_sel & vns_videooverlaysoc_interface0_bank_bus_we) & (vns_videooverlaysoc_interface0_bank_bus_adr[3:0] == 3'd7));
assign vns_videooverlaysoc_csrbank0_bus_errors0_r = vns_videooverlaysoc_interface0_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank0_bus_errors0_re = ((vns_videooverlaysoc_csrbank0_sel & vns_videooverlaysoc_interface0_bank_bus_we) & (vns_videooverlaysoc_interface0_bank_bus_adr[3:0] == 4'd8));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full[31:0];
assign vns_videooverlaysoc_csrbank0_scratch3_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full[31:24];
assign vns_videooverlaysoc_csrbank0_scratch2_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full[23:16];
assign vns_videooverlaysoc_csrbank0_scratch1_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full[15:8];
assign vns_videooverlaysoc_csrbank0_scratch0_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full[7:0];
assign vns_videooverlaysoc_csrbank0_bus_errors3_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors_status[31:24];
assign vns_videooverlaysoc_csrbank0_bus_errors2_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors_status[23:16];
assign vns_videooverlaysoc_csrbank0_bus_errors1_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors_status[15:8];
assign vns_videooverlaysoc_csrbank0_bus_errors0_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors_status[7:0];
assign vns_videooverlaysoc_csrbank1_sel = (vns_videooverlaysoc_interface1_bank_bus_adr[13:9] == 4'd10);
assign vns_videooverlaysoc_csrbank1_half_sys8x_taps0_r = vns_videooverlaysoc_interface1_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank1_half_sys8x_taps0_re = ((vns_videooverlaysoc_csrbank1_sel & vns_videooverlaysoc_interface1_bank_bus_we) & (vns_videooverlaysoc_interface1_bank_bus_adr[2:0] == 1'd0));
assign vns_videooverlaysoc_csrbank1_dly_sel0_r = vns_videooverlaysoc_interface1_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank1_dly_sel0_re = ((vns_videooverlaysoc_csrbank1_sel & vns_videooverlaysoc_interface1_bank_bus_we) & (vns_videooverlaysoc_interface1_bank_bus_adr[2:0] == 1'd1));
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_r = vns_videooverlaysoc_interface1_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re = ((vns_videooverlaysoc_csrbank1_sel & vns_videooverlaysoc_interface1_bank_bus_we) & (vns_videooverlaysoc_interface1_bank_bus_adr[2:0] == 2'd2));
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_r = vns_videooverlaysoc_interface1_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re = ((vns_videooverlaysoc_csrbank1_sel & vns_videooverlaysoc_interface1_bank_bus_we) & (vns_videooverlaysoc_interface1_bank_bus_adr[2:0] == 2'd3));
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_r = vns_videooverlaysoc_interface1_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re = ((vns_videooverlaysoc_csrbank1_sel & vns_videooverlaysoc_interface1_bank_bus_we) & (vns_videooverlaysoc_interface1_bank_bus_adr[2:0] == 3'd4));
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_r = vns_videooverlaysoc_interface1_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re = ((vns_videooverlaysoc_csrbank1_sel & vns_videooverlaysoc_interface1_bank_bus_we) & (vns_videooverlaysoc_interface1_bank_bus_adr[2:0] == 3'd5));
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_half_sys8x_taps_storage = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_half_sys8x_taps_storage_full[3:0];
assign vns_videooverlaysoc_csrbank1_half_sys8x_taps0_w = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_half_sys8x_taps_storage_full[3:0];
assign soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage_full[3:0];
assign vns_videooverlaysoc_csrbank1_dly_sel0_w = soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage_full[3:0];
assign vns_videooverlaysoc_csrbank2_sel = (vns_videooverlaysoc_interface2_bank_bus_adr[13:9] == 5'd21);
assign vns_videooverlaysoc_csrbank2_Km6_r = vns_videooverlaysoc_interface2_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank2_Km6_re = ((vns_videooverlaysoc_csrbank2_sel & vns_videooverlaysoc_interface2_bank_bus_we) & (vns_videooverlaysoc_interface2_bank_bus_adr[3:0] == 1'd0));
assign vns_videooverlaysoc_csrbank2_Km5_r = vns_videooverlaysoc_interface2_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank2_Km5_re = ((vns_videooverlaysoc_csrbank2_sel & vns_videooverlaysoc_interface2_bank_bus_we) & (vns_videooverlaysoc_interface2_bank_bus_adr[3:0] == 1'd1));
assign vns_videooverlaysoc_csrbank2_Km4_r = vns_videooverlaysoc_interface2_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank2_Km4_re = ((vns_videooverlaysoc_csrbank2_sel & vns_videooverlaysoc_interface2_bank_bus_we) & (vns_videooverlaysoc_interface2_bank_bus_adr[3:0] == 2'd2));
assign vns_videooverlaysoc_csrbank2_Km3_r = vns_videooverlaysoc_interface2_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank2_Km3_re = ((vns_videooverlaysoc_csrbank2_sel & vns_videooverlaysoc_interface2_bank_bus_we) & (vns_videooverlaysoc_interface2_bank_bus_adr[3:0] == 2'd3));
assign vns_videooverlaysoc_csrbank2_Km2_r = vns_videooverlaysoc_interface2_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank2_Km2_re = ((vns_videooverlaysoc_csrbank2_sel & vns_videooverlaysoc_interface2_bank_bus_we) & (vns_videooverlaysoc_interface2_bank_bus_adr[3:0] == 3'd4));
assign vns_videooverlaysoc_csrbank2_Km1_r = vns_videooverlaysoc_interface2_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank2_Km1_re = ((vns_videooverlaysoc_csrbank2_sel & vns_videooverlaysoc_interface2_bank_bus_we) & (vns_videooverlaysoc_interface2_bank_bus_adr[3:0] == 3'd5));
assign vns_videooverlaysoc_csrbank2_Km0_r = vns_videooverlaysoc_interface2_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank2_Km0_re = ((vns_videooverlaysoc_csrbank2_sel & vns_videooverlaysoc_interface2_bank_bus_we) & (vns_videooverlaysoc_interface2_bank_bus_adr[3:0] == 3'd6));
assign vns_videooverlaysoc_csrbank2_Km_valid0_r = vns_videooverlaysoc_interface2_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank2_Km_valid0_re = ((vns_videooverlaysoc_csrbank2_sel & vns_videooverlaysoc_interface2_bank_bus_we) & (vns_videooverlaysoc_interface2_bank_bus_adr[3:0] == 3'd7));
assign vns_videooverlaysoc_csrbank2_hpd_ena0_r = vns_videooverlaysoc_interface2_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank2_hpd_ena0_re = ((vns_videooverlaysoc_csrbank2_sel & vns_videooverlaysoc_interface2_bank_bus_we) & (vns_videooverlaysoc_interface2_bank_bus_adr[3:0] == 4'd8));
assign soc_videooverlaysoc_hdcp_Km_storage = soc_videooverlaysoc_hdcp_Km_storage_full[55:0];
assign vns_videooverlaysoc_csrbank2_Km6_w = soc_videooverlaysoc_hdcp_Km_storage_full[55:48];
assign vns_videooverlaysoc_csrbank2_Km5_w = soc_videooverlaysoc_hdcp_Km_storage_full[47:40];
assign vns_videooverlaysoc_csrbank2_Km4_w = soc_videooverlaysoc_hdcp_Km_storage_full[39:32];
assign vns_videooverlaysoc_csrbank2_Km3_w = soc_videooverlaysoc_hdcp_Km_storage_full[31:24];
assign vns_videooverlaysoc_csrbank2_Km2_w = soc_videooverlaysoc_hdcp_Km_storage_full[23:16];
assign vns_videooverlaysoc_csrbank2_Km1_w = soc_videooverlaysoc_hdcp_Km_storage_full[15:8];
assign vns_videooverlaysoc_csrbank2_Km0_w = soc_videooverlaysoc_hdcp_Km_storage_full[7:0];
assign soc_videooverlaysoc_hdcp_Km_valid_storage = soc_videooverlaysoc_hdcp_Km_valid_storage_full;
assign vns_videooverlaysoc_csrbank2_Km_valid0_w = soc_videooverlaysoc_hdcp_Km_valid_storage_full;
assign soc_videooverlaysoc_hdcp_hpd_ena_storage = soc_videooverlaysoc_hdcp_hpd_ena_storage_full;
assign vns_videooverlaysoc_csrbank2_hpd_ena0_w = soc_videooverlaysoc_hdcp_hpd_ena_storage_full;
assign vns_videooverlaysoc_csrbank3_sel = (vns_videooverlaysoc_interface3_bank_bus_adr[13:9] == 4'd13);
assign vns_videooverlaysoc_csrbank3_underflow_enable0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank3_underflow_enable0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 1'd0));
assign soc_videooverlaysoc_hdmi_core_out0_underflow_update_underflow_update_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_core_out0_underflow_update_underflow_update_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 1'd1));
assign vns_videooverlaysoc_csrbank3_underflow_counter3_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_underflow_counter3_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 2'd2));
assign vns_videooverlaysoc_csrbank3_underflow_counter2_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_underflow_counter2_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 2'd3));
assign vns_videooverlaysoc_csrbank3_underflow_counter1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_underflow_counter1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 3'd4));
assign vns_videooverlaysoc_csrbank3_underflow_counter0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_underflow_counter0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 3'd5));
assign vns_videooverlaysoc_csrbank3_initiator_enable0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank3_initiator_enable0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 3'd6));
assign vns_videooverlaysoc_csrbank3_initiator_hres1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank3_initiator_hres1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 3'd7));
assign vns_videooverlaysoc_csrbank3_initiator_hres0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_hres0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 4'd8));
assign vns_videooverlaysoc_csrbank3_initiator_hsync_start1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank3_initiator_hsync_start1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 4'd9));
assign vns_videooverlaysoc_csrbank3_initiator_hsync_start0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_hsync_start0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 4'd10));
assign vns_videooverlaysoc_csrbank3_initiator_hsync_end1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank3_initiator_hsync_end1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 4'd11));
assign vns_videooverlaysoc_csrbank3_initiator_hsync_end0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_hsync_end0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 4'd12));
assign vns_videooverlaysoc_csrbank3_initiator_hscan1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank3_initiator_hscan1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 4'd13));
assign vns_videooverlaysoc_csrbank3_initiator_hscan0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_hscan0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 4'd14));
assign vns_videooverlaysoc_csrbank3_initiator_vres1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank3_initiator_vres1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 4'd15));
assign vns_videooverlaysoc_csrbank3_initiator_vres0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_vres0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd16));
assign vns_videooverlaysoc_csrbank3_initiator_vsync_start1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank3_initiator_vsync_start1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd17));
assign vns_videooverlaysoc_csrbank3_initiator_vsync_start0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_vsync_start0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd18));
assign vns_videooverlaysoc_csrbank3_initiator_vsync_end1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank3_initiator_vsync_end1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd19));
assign vns_videooverlaysoc_csrbank3_initiator_vsync_end0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_vsync_end0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd20));
assign vns_videooverlaysoc_csrbank3_initiator_vscan1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank3_initiator_vscan1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd21));
assign vns_videooverlaysoc_csrbank3_initiator_vscan0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_vscan0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd22));
assign vns_videooverlaysoc_csrbank3_initiator_base3_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_base3_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd23));
assign vns_videooverlaysoc_csrbank3_initiator_base2_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_base2_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd24));
assign vns_videooverlaysoc_csrbank3_initiator_base1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_base1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd25));
assign vns_videooverlaysoc_csrbank3_initiator_base0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_base0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd26));
assign vns_videooverlaysoc_csrbank3_initiator_length3_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_length3_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd27));
assign vns_videooverlaysoc_csrbank3_initiator_length2_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_length2_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd28));
assign vns_videooverlaysoc_csrbank3_initiator_length1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_length1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd29));
assign vns_videooverlaysoc_csrbank3_initiator_length0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_initiator_length0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd30));
assign vns_videooverlaysoc_csrbank3_dma_delay_base3_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_dma_delay_base3_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 5'd31));
assign vns_videooverlaysoc_csrbank3_dma_delay_base2_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_dma_delay_base2_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 6'd32));
assign vns_videooverlaysoc_csrbank3_dma_delay_base1_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_dma_delay_base1_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 6'd33));
assign vns_videooverlaysoc_csrbank3_dma_delay_base0_r = vns_videooverlaysoc_interface3_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank3_dma_delay_base0_re = ((vns_videooverlaysoc_csrbank3_sel & vns_videooverlaysoc_interface3_bank_bus_we) & (vns_videooverlaysoc_interface3_bank_bus_adr[5:0] == 6'd34));
assign soc_videooverlaysoc_hdmi_core_out0_underflow_enable_storage = soc_videooverlaysoc_hdmi_core_out0_underflow_enable_storage_full;
assign vns_videooverlaysoc_csrbank3_underflow_enable0_w = soc_videooverlaysoc_hdmi_core_out0_underflow_enable_storage_full;
assign vns_videooverlaysoc_csrbank3_underflow_counter3_w = soc_videooverlaysoc_hdmi_core_out0_underflow_counter_status[31:24];
assign vns_videooverlaysoc_csrbank3_underflow_counter2_w = soc_videooverlaysoc_hdmi_core_out0_underflow_counter_status[23:16];
assign vns_videooverlaysoc_csrbank3_underflow_counter1_w = soc_videooverlaysoc_hdmi_core_out0_underflow_counter_status[15:8];
assign vns_videooverlaysoc_csrbank3_underflow_counter0_w = soc_videooverlaysoc_hdmi_core_out0_underflow_counter_status[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_enable_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_enable_storage_full;
assign vns_videooverlaysoc_csrbank3_initiator_enable0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_enable_storage_full;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_storage_full[11:0];
assign vns_videooverlaysoc_csrbank3_initiator_hres1_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_storage_full[11:8];
assign vns_videooverlaysoc_csrbank3_initiator_hres0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_storage_full[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_storage_full[11:0];
assign vns_videooverlaysoc_csrbank3_initiator_hsync_start1_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_storage_full[11:8];
assign vns_videooverlaysoc_csrbank3_initiator_hsync_start0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_storage_full[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_storage_full[11:0];
assign vns_videooverlaysoc_csrbank3_initiator_hsync_end1_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_storage_full[11:8];
assign vns_videooverlaysoc_csrbank3_initiator_hsync_end0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_storage_full[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_storage_full[11:0];
assign vns_videooverlaysoc_csrbank3_initiator_hscan1_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_storage_full[11:8];
assign vns_videooverlaysoc_csrbank3_initiator_hscan0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_storage_full[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_storage_full[11:0];
assign vns_videooverlaysoc_csrbank3_initiator_vres1_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_storage_full[11:8];
assign vns_videooverlaysoc_csrbank3_initiator_vres0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_storage_full[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_storage_full[11:0];
assign vns_videooverlaysoc_csrbank3_initiator_vsync_start1_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_storage_full[11:8];
assign vns_videooverlaysoc_csrbank3_initiator_vsync_start0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_storage_full[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_storage_full[11:0];
assign vns_videooverlaysoc_csrbank3_initiator_vsync_end1_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_storage_full[11:8];
assign vns_videooverlaysoc_csrbank3_initiator_vsync_end0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_storage_full[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_storage_full[11:0];
assign vns_videooverlaysoc_csrbank3_initiator_vscan1_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_storage_full[11:8];
assign vns_videooverlaysoc_csrbank3_initiator_vscan0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_storage_full[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage_full[31:0];
assign vns_videooverlaysoc_csrbank3_initiator_base3_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage_full[31:24];
assign vns_videooverlaysoc_csrbank3_initiator_base2_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage_full[23:16];
assign vns_videooverlaysoc_csrbank3_initiator_base1_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage_full[15:8];
assign vns_videooverlaysoc_csrbank3_initiator_base0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage_full[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage_full[31:0];
assign vns_videooverlaysoc_csrbank3_initiator_length3_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage_full[31:24];
assign vns_videooverlaysoc_csrbank3_initiator_length2_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage_full[23:16];
assign vns_videooverlaysoc_csrbank3_initiator_length1_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage_full[15:8];
assign vns_videooverlaysoc_csrbank3_initiator_length0_w = soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage_full[7:0];
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_storage = soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full[31:0];
assign vns_videooverlaysoc_csrbank3_dma_delay_base3_w = soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full[31:24];
assign vns_videooverlaysoc_csrbank3_dma_delay_base2_w = soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full[23:16];
assign vns_videooverlaysoc_csrbank3_dma_delay_base1_w = soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full[15:8];
assign vns_videooverlaysoc_csrbank3_dma_delay_base0_w = soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full[7:0];
assign vns_videooverlaysoc_sram0_sel = (vns_videooverlaysoc_interface0_sram_bus_adr[13:9] == 5'd16);
always @(*) begin
	vns_videooverlaysoc_interface0_sram_bus_dat_r <= 8'd0;
	if (vns_videooverlaysoc_sram0_sel_r) begin
		vns_videooverlaysoc_interface0_sram_bus_dat_r <= vns_videooverlaysoc_sram0_dat_r;
	end
end
assign vns_videooverlaysoc_sram0_we = (vns_videooverlaysoc_sram0_sel & vns_videooverlaysoc_interface0_sram_bus_we);
assign vns_videooverlaysoc_sram0_dat_w = vns_videooverlaysoc_interface0_sram_bus_dat_w;
assign vns_videooverlaysoc_sram0_adr = vns_videooverlaysoc_interface0_sram_bus_adr[7:0];
assign vns_videooverlaysoc_csrbank4_sel = (vns_videooverlaysoc_interface4_bank_bus_adr[13:9] == 4'd14);
assign vns_videooverlaysoc_csrbank4_edid_hpd_notif_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_edid_hpd_notif_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 1'd0));
assign vns_videooverlaysoc_csrbank4_edid_hpd_en0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_edid_hpd_en0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 1'd1));
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_reset0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_reset0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 2'd2));
assign vns_videooverlaysoc_csrbank4_clocking_locked_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_clocking_locked_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 2'd3));
assign soc_videooverlaysoc_hdmi_in0_mmcm_read_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in0_mmcm_read_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 3'd4));
assign soc_videooverlaysoc_hdmi_in0_mmcm_write_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in0_mmcm_write_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 3'd5));
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 3'd6));
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_adr0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[6:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_adr0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 3'd7));
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w1_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w1_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 4'd8));
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 4'd9));
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r1_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r1_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 4'd10));
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 4'd11));
assign soc_videooverlaysoc_hdmi_in0_mmcm_write_o_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in0_mmcm_write_o_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 4'd12));
assign soc_videooverlaysoc_hdmi_in0_mmcm_read_o_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in0_mmcm_read_o_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 4'd13));
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r1_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r1_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 4'd14));
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 4'd15));
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_o_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_o_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd16));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[4:0];
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd17));
assign vns_videooverlaysoc_csrbank4_data0_cap_phase_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[1:0];
assign vns_videooverlaysoc_csrbank4_data0_cap_phase_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd18));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_phase_reset_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_phase_reset_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd19));
assign vns_videooverlaysoc_csrbank4_data0_charsync_char_synced_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_data0_charsync_char_synced_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd20));
assign vns_videooverlaysoc_csrbank4_data0_charsync_ctl_pos_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank4_data0_charsync_ctl_pos_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd21));
assign soc_videooverlaysoc_hdmi_in0_wer0_update_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in0_wer0_update_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd22));
assign vns_videooverlaysoc_csrbank4_data0_wer_value2_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_data0_wer_value2_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd23));
assign vns_videooverlaysoc_csrbank4_data0_wer_value1_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_data0_wer_value1_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd24));
assign vns_videooverlaysoc_csrbank4_data0_wer_value0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_data0_wer_value0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd25));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[4:0];
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd26));
assign vns_videooverlaysoc_csrbank4_data1_cap_phase_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[1:0];
assign vns_videooverlaysoc_csrbank4_data1_cap_phase_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd27));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_phase_reset_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_phase_reset_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd28));
assign vns_videooverlaysoc_csrbank4_data1_charsync_char_synced_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_data1_charsync_char_synced_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd29));
assign vns_videooverlaysoc_csrbank4_data1_charsync_ctl_pos_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank4_data1_charsync_ctl_pos_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd30));
assign soc_videooverlaysoc_hdmi_in0_wer1_update_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in0_wer1_update_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 5'd31));
assign vns_videooverlaysoc_csrbank4_data1_wer_value2_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_data1_wer_value2_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd32));
assign vns_videooverlaysoc_csrbank4_data1_wer_value1_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_data1_wer_value1_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd33));
assign vns_videooverlaysoc_csrbank4_data1_wer_value0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_data1_wer_value0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd34));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[4:0];
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd35));
assign vns_videooverlaysoc_csrbank4_data2_cap_phase_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[1:0];
assign vns_videooverlaysoc_csrbank4_data2_cap_phase_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd36));
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_phase_reset_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_phase_reset_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd37));
assign vns_videooverlaysoc_csrbank4_data2_charsync_char_synced_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_data2_charsync_char_synced_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd38));
assign vns_videooverlaysoc_csrbank4_data2_charsync_ctl_pos_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank4_data2_charsync_ctl_pos_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd39));
assign soc_videooverlaysoc_hdmi_in0_wer2_update_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in0_wer2_update_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd40));
assign vns_videooverlaysoc_csrbank4_data2_wer_value2_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_data2_wer_value2_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd41));
assign vns_videooverlaysoc_csrbank4_data2_wer_value1_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_data2_wer_value1_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd42));
assign vns_videooverlaysoc_csrbank4_data2_wer_value0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_data2_wer_value0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd43));
assign vns_videooverlaysoc_csrbank4_chansync_channels_synced_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_chansync_channels_synced_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd44));
assign vns_videooverlaysoc_csrbank4_decode_terc4_dvimode0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank4_decode_terc4_dvimode0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd45));
assign vns_videooverlaysoc_csrbank4_resdetection_hres1_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[2:0];
assign vns_videooverlaysoc_csrbank4_resdetection_hres1_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd46));
assign vns_videooverlaysoc_csrbank4_resdetection_hres0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_resdetection_hres0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd47));
assign vns_videooverlaysoc_csrbank4_resdetection_vres1_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[2:0];
assign vns_videooverlaysoc_csrbank4_resdetection_vres1_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd48));
assign vns_videooverlaysoc_csrbank4_resdetection_vres0_r = vns_videooverlaysoc_interface4_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank4_resdetection_vres0_re = ((vns_videooverlaysoc_csrbank4_sel & vns_videooverlaysoc_interface4_bank_bus_we) & (vns_videooverlaysoc_interface4_bank_bus_adr[5:0] == 6'd49));
assign vns_videooverlaysoc_csrbank4_edid_hpd_notif_w = soc_videooverlaysoc_hdmi_in0_edid_status;
assign soc_videooverlaysoc_hdmi_in0_edid_storage = soc_videooverlaysoc_hdmi_in0_edid_storage_full;
assign vns_videooverlaysoc_csrbank4_edid_hpd_en0_w = soc_videooverlaysoc_hdmi_in0_edid_storage_full;
assign soc_videooverlaysoc_hdmi_in0_mmcm_reset_storage = soc_videooverlaysoc_hdmi_in0_mmcm_reset_storage_full;
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_reset0_w = soc_videooverlaysoc_hdmi_in0_mmcm_reset_storage_full;
assign vns_videooverlaysoc_csrbank4_clocking_locked_w = soc_videooverlaysoc_hdmi_in0_locked_status;
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_w = soc_videooverlaysoc_hdmi_in0_mmcm_drdy_status;
assign soc_videooverlaysoc_hdmi_in0_mmcm_adr_storage = soc_videooverlaysoc_hdmi_in0_mmcm_adr_storage_full[6:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_adr0_w = soc_videooverlaysoc_hdmi_in0_mmcm_adr_storage_full[6:0];
assign soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage = soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage_full[15:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w1_w = soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage_full[15:8];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w0_w = soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage_full[7:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r1_w = soc_videooverlaysoc_hdmi_in0_mmcm_dat_r_status[15:8];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r0_w = soc_videooverlaysoc_hdmi_in0_mmcm_dat_r_status[7:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r1_w = soc_videooverlaysoc_hdmi_in0_mmcm_dat_o_r_status[15:8];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r0_w = soc_videooverlaysoc_hdmi_in0_mmcm_dat_o_r_status[7:0];
assign vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_o_w = soc_videooverlaysoc_hdmi_in0_mmcm_drdy_o_status;
assign vns_videooverlaysoc_csrbank4_data0_cap_phase_w = soc_videooverlaysoc_hdmi_in0_s7datacapture0_status[1:0];
assign vns_videooverlaysoc_csrbank4_data0_charsync_char_synced_w = soc_videooverlaysoc_hdmi_in0_charsync0_char_synced_status;
assign vns_videooverlaysoc_csrbank4_data0_charsync_ctl_pos_w = soc_videooverlaysoc_hdmi_in0_charsync0_ctl_pos_status[3:0];
assign vns_videooverlaysoc_csrbank4_data0_wer_value2_w = soc_videooverlaysoc_hdmi_in0_wer0_status[23:16];
assign vns_videooverlaysoc_csrbank4_data0_wer_value1_w = soc_videooverlaysoc_hdmi_in0_wer0_status[15:8];
assign vns_videooverlaysoc_csrbank4_data0_wer_value0_w = soc_videooverlaysoc_hdmi_in0_wer0_status[7:0];
assign vns_videooverlaysoc_csrbank4_data1_cap_phase_w = soc_videooverlaysoc_hdmi_in0_s7datacapture1_status[1:0];
assign vns_videooverlaysoc_csrbank4_data1_charsync_char_synced_w = soc_videooverlaysoc_hdmi_in0_charsync1_char_synced_status;
assign vns_videooverlaysoc_csrbank4_data1_charsync_ctl_pos_w = soc_videooverlaysoc_hdmi_in0_charsync1_ctl_pos_status[3:0];
assign vns_videooverlaysoc_csrbank4_data1_wer_value2_w = soc_videooverlaysoc_hdmi_in0_wer1_status[23:16];
assign vns_videooverlaysoc_csrbank4_data1_wer_value1_w = soc_videooverlaysoc_hdmi_in0_wer1_status[15:8];
assign vns_videooverlaysoc_csrbank4_data1_wer_value0_w = soc_videooverlaysoc_hdmi_in0_wer1_status[7:0];
assign vns_videooverlaysoc_csrbank4_data2_cap_phase_w = soc_videooverlaysoc_hdmi_in0_s7datacapture2_status[1:0];
assign vns_videooverlaysoc_csrbank4_data2_charsync_char_synced_w = soc_videooverlaysoc_hdmi_in0_charsync2_char_synced_status;
assign vns_videooverlaysoc_csrbank4_data2_charsync_ctl_pos_w = soc_videooverlaysoc_hdmi_in0_charsync2_ctl_pos_status[3:0];
assign vns_videooverlaysoc_csrbank4_data2_wer_value2_w = soc_videooverlaysoc_hdmi_in0_wer2_status[23:16];
assign vns_videooverlaysoc_csrbank4_data2_wer_value1_w = soc_videooverlaysoc_hdmi_in0_wer2_status[15:8];
assign vns_videooverlaysoc_csrbank4_data2_wer_value0_w = soc_videooverlaysoc_hdmi_in0_wer2_status[7:0];
assign vns_videooverlaysoc_csrbank4_chansync_channels_synced_w = soc_videooverlaysoc_hdmi_in0_chansync_status;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_storage = soc_videooverlaysoc_hdmi_in0_decode_terc4_storage_full;
assign vns_videooverlaysoc_csrbank4_decode_terc4_dvimode0_w = soc_videooverlaysoc_hdmi_in0_decode_terc4_storage_full;
assign vns_videooverlaysoc_csrbank4_resdetection_hres1_w = soc_videooverlaysoc_hdmi_in0_resdetection_hres_status[10:8];
assign vns_videooverlaysoc_csrbank4_resdetection_hres0_w = soc_videooverlaysoc_hdmi_in0_resdetection_hres_status[7:0];
assign vns_videooverlaysoc_csrbank4_resdetection_vres1_w = soc_videooverlaysoc_hdmi_in0_resdetection_vres_status[10:8];
assign vns_videooverlaysoc_csrbank4_resdetection_vres0_w = soc_videooverlaysoc_hdmi_in0_resdetection_vres_status[7:0];
assign vns_videooverlaysoc_csrbank5_sel = (vns_videooverlaysoc_interface5_bank_bus_adr[13:9] == 4'd15);
assign vns_videooverlaysoc_csrbank5_value3_r = vns_videooverlaysoc_interface5_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank5_value3_re = ((vns_videooverlaysoc_csrbank5_sel & vns_videooverlaysoc_interface5_bank_bus_we) & (vns_videooverlaysoc_interface5_bank_bus_adr[1:0] == 1'd0));
assign vns_videooverlaysoc_csrbank5_value2_r = vns_videooverlaysoc_interface5_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank5_value2_re = ((vns_videooverlaysoc_csrbank5_sel & vns_videooverlaysoc_interface5_bank_bus_we) & (vns_videooverlaysoc_interface5_bank_bus_adr[1:0] == 1'd1));
assign vns_videooverlaysoc_csrbank5_value1_r = vns_videooverlaysoc_interface5_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank5_value1_re = ((vns_videooverlaysoc_csrbank5_sel & vns_videooverlaysoc_interface5_bank_bus_we) & (vns_videooverlaysoc_interface5_bank_bus_adr[1:0] == 2'd2));
assign vns_videooverlaysoc_csrbank5_value0_r = vns_videooverlaysoc_interface5_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank5_value0_re = ((vns_videooverlaysoc_csrbank5_sel & vns_videooverlaysoc_interface5_bank_bus_we) & (vns_videooverlaysoc_interface5_bank_bus_adr[1:0] == 2'd3));
assign vns_videooverlaysoc_csrbank5_value3_w = soc_videooverlaysoc_hdmi_in0_freq_status[31:24];
assign vns_videooverlaysoc_csrbank5_value2_w = soc_videooverlaysoc_hdmi_in0_freq_status[23:16];
assign vns_videooverlaysoc_csrbank5_value1_w = soc_videooverlaysoc_hdmi_in0_freq_status[15:8];
assign vns_videooverlaysoc_csrbank5_value0_w = soc_videooverlaysoc_hdmi_in0_freq_status[7:0];
assign vns_videooverlaysoc_sram1_sel = (vns_videooverlaysoc_interface1_sram_bus_adr[13:9] == 5'd19);
always @(*) begin
	vns_videooverlaysoc_interface1_sram_bus_dat_r <= 8'd0;
	if (vns_videooverlaysoc_sram1_sel_r) begin
		vns_videooverlaysoc_interface1_sram_bus_dat_r <= vns_videooverlaysoc_sram1_dat_r;
	end
end
assign vns_videooverlaysoc_sram1_we = (vns_videooverlaysoc_sram1_sel & vns_videooverlaysoc_interface1_sram_bus_we);
assign vns_videooverlaysoc_sram1_dat_w = vns_videooverlaysoc_interface1_sram_bus_dat_w;
assign vns_videooverlaysoc_sram1_adr = vns_videooverlaysoc_interface1_sram_bus_adr[7:0];
assign vns_videooverlaysoc_csrbank6_sel = (vns_videooverlaysoc_interface6_bank_bus_adr[13:9] == 5'd17);
assign vns_videooverlaysoc_csrbank6_edid_hpd_notif_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank6_edid_hpd_notif_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 1'd0));
assign vns_videooverlaysoc_csrbank6_edid_hpd_en0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank6_edid_hpd_en0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 1'd1));
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_reset0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_reset0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 2'd2));
assign vns_videooverlaysoc_csrbank6_clocking_locked_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank6_clocking_locked_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 2'd3));
assign soc_videooverlaysoc_hdmi_in1_mmcm_read_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in1_mmcm_read_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 3'd4));
assign soc_videooverlaysoc_hdmi_in1_mmcm_write_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in1_mmcm_write_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 3'd5));
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_drdy_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_drdy_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 3'd6));
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_adr0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[6:0];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_adr0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 3'd7));
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w1_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w1_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 4'd8));
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 4'd9));
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r1_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r1_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 4'd10));
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 4'd11));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[4:0];
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 4'd12));
assign vns_videooverlaysoc_csrbank6_data0_cap_phase_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[1:0];
assign vns_videooverlaysoc_csrbank6_data0_cap_phase_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 4'd13));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_phase_reset_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_phase_reset_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 4'd14));
assign vns_videooverlaysoc_csrbank6_data0_charsync_char_synced_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank6_data0_charsync_char_synced_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 4'd15));
assign vns_videooverlaysoc_csrbank6_data0_charsync_ctl_pos_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank6_data0_charsync_ctl_pos_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd16));
assign soc_videooverlaysoc_hdmi_in1_wer0_update_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in1_wer0_update_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd17));
assign vns_videooverlaysoc_csrbank6_data0_wer_value2_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_data0_wer_value2_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd18));
assign vns_videooverlaysoc_csrbank6_data0_wer_value1_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_data0_wer_value1_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd19));
assign vns_videooverlaysoc_csrbank6_data0_wer_value0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_data0_wer_value0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd20));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[4:0];
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd21));
assign vns_videooverlaysoc_csrbank6_data1_cap_phase_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[1:0];
assign vns_videooverlaysoc_csrbank6_data1_cap_phase_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd22));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_phase_reset_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_phase_reset_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd23));
assign vns_videooverlaysoc_csrbank6_data1_charsync_char_synced_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank6_data1_charsync_char_synced_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd24));
assign vns_videooverlaysoc_csrbank6_data1_charsync_ctl_pos_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank6_data1_charsync_ctl_pos_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd25));
assign soc_videooverlaysoc_hdmi_in1_wer1_update_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in1_wer1_update_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd26));
assign vns_videooverlaysoc_csrbank6_data1_wer_value2_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_data1_wer_value2_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd27));
assign vns_videooverlaysoc_csrbank6_data1_wer_value1_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_data1_wer_value1_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd28));
assign vns_videooverlaysoc_csrbank6_data1_wer_value0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_data1_wer_value0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd29));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[4:0];
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd30));
assign vns_videooverlaysoc_csrbank6_data2_cap_phase_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[1:0];
assign vns_videooverlaysoc_csrbank6_data2_cap_phase_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 5'd31));
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_phase_reset_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_phase_reset_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd32));
assign vns_videooverlaysoc_csrbank6_data2_charsync_char_synced_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank6_data2_charsync_char_synced_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd33));
assign vns_videooverlaysoc_csrbank6_data2_charsync_ctl_pos_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank6_data2_charsync_ctl_pos_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd34));
assign soc_videooverlaysoc_hdmi_in1_wer2_update_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in1_wer2_update_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd35));
assign vns_videooverlaysoc_csrbank6_data2_wer_value2_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_data2_wer_value2_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd36));
assign vns_videooverlaysoc_csrbank6_data2_wer_value1_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_data2_wer_value1_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd37));
assign vns_videooverlaysoc_csrbank6_data2_wer_value0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_data2_wer_value0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd38));
assign vns_videooverlaysoc_csrbank6_chansync_channels_synced_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank6_chansync_channels_synced_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd39));
assign vns_videooverlaysoc_csrbank6_decode_terc4_dvimode0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank6_decode_terc4_dvimode0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd40));
assign vns_videooverlaysoc_csrbank6_resdetection_hres1_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[2:0];
assign vns_videooverlaysoc_csrbank6_resdetection_hres1_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd41));
assign vns_videooverlaysoc_csrbank6_resdetection_hres0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_resdetection_hres0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd42));
assign vns_videooverlaysoc_csrbank6_resdetection_vres1_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[2:0];
assign vns_videooverlaysoc_csrbank6_resdetection_vres1_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd43));
assign vns_videooverlaysoc_csrbank6_resdetection_vres0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_resdetection_vres0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd44));
assign soc_videooverlaysoc_hdmi_in1_frame_overflow_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[0];
assign soc_videooverlaysoc_hdmi_in1_frame_overflow_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd45));
assign vns_videooverlaysoc_csrbank6_dma_frame_size3_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[4:0];
assign vns_videooverlaysoc_csrbank6_dma_frame_size3_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd46));
assign vns_videooverlaysoc_csrbank6_dma_frame_size2_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_dma_frame_size2_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd47));
assign vns_videooverlaysoc_csrbank6_dma_frame_size1_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_dma_frame_size1_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd48));
assign vns_videooverlaysoc_csrbank6_dma_frame_size0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_dma_frame_size0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd49));
assign vns_videooverlaysoc_csrbank6_dma_slot0_status0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[1:0];
assign vns_videooverlaysoc_csrbank6_dma_slot0_status0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd50));
assign vns_videooverlaysoc_csrbank6_dma_slot0_address3_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[4:0];
assign vns_videooverlaysoc_csrbank6_dma_slot0_address3_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd51));
assign vns_videooverlaysoc_csrbank6_dma_slot0_address2_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_dma_slot0_address2_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd52));
assign vns_videooverlaysoc_csrbank6_dma_slot0_address1_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_dma_slot0_address1_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd53));
assign vns_videooverlaysoc_csrbank6_dma_slot0_address0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_dma_slot0_address0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd54));
assign vns_videooverlaysoc_csrbank6_dma_slot1_status0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[1:0];
assign vns_videooverlaysoc_csrbank6_dma_slot1_status0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd55));
assign vns_videooverlaysoc_csrbank6_dma_slot1_address3_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[4:0];
assign vns_videooverlaysoc_csrbank6_dma_slot1_address3_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd56));
assign vns_videooverlaysoc_csrbank6_dma_slot1_address2_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_dma_slot1_address2_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd57));
assign vns_videooverlaysoc_csrbank6_dma_slot1_address1_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_dma_slot1_address1_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd58));
assign vns_videooverlaysoc_csrbank6_dma_slot1_address0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank6_dma_slot1_address0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd59));
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_status_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[1:0];
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_status_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd60));
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[1:0];
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd61));
assign vns_videooverlaysoc_csrbank6_dma_ev_enable0_r = vns_videooverlaysoc_interface6_bank_bus_dat_w[1:0];
assign vns_videooverlaysoc_csrbank6_dma_ev_enable0_re = ((vns_videooverlaysoc_csrbank6_sel & vns_videooverlaysoc_interface6_bank_bus_we) & (vns_videooverlaysoc_interface6_bank_bus_adr[5:0] == 6'd62));
assign vns_videooverlaysoc_csrbank6_edid_hpd_notif_w = soc_videooverlaysoc_hdmi_in1_edid_status;
assign soc_videooverlaysoc_hdmi_in1_edid_storage = soc_videooverlaysoc_hdmi_in1_edid_storage_full;
assign vns_videooverlaysoc_csrbank6_edid_hpd_en0_w = soc_videooverlaysoc_hdmi_in1_edid_storage_full;
assign soc_videooverlaysoc_hdmi_in1_mmcm_reset_storage = soc_videooverlaysoc_hdmi_in1_mmcm_reset_storage_full;
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_reset0_w = soc_videooverlaysoc_hdmi_in1_mmcm_reset_storage_full;
assign vns_videooverlaysoc_csrbank6_clocking_locked_w = soc_videooverlaysoc_hdmi_in1_locked_status;
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_drdy_w = soc_videooverlaysoc_hdmi_in1_mmcm_drdy_status;
assign soc_videooverlaysoc_hdmi_in1_mmcm_adr_storage = soc_videooverlaysoc_hdmi_in1_mmcm_adr_storage_full[6:0];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_adr0_w = soc_videooverlaysoc_hdmi_in1_mmcm_adr_storage_full[6:0];
assign soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_storage = soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_storage_full[15:0];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w1_w = soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_storage_full[15:8];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w0_w = soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_storage_full[7:0];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r1_w = soc_videooverlaysoc_hdmi_in1_mmcm_dat_r_status[15:8];
assign vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r0_w = soc_videooverlaysoc_hdmi_in1_mmcm_dat_r_status[7:0];
assign vns_videooverlaysoc_csrbank6_data0_cap_phase_w = soc_videooverlaysoc_hdmi_in1_s7datacapture0_status[1:0];
assign vns_videooverlaysoc_csrbank6_data0_charsync_char_synced_w = soc_videooverlaysoc_hdmi_in1_charsync0_char_synced_status;
assign vns_videooverlaysoc_csrbank6_data0_charsync_ctl_pos_w = soc_videooverlaysoc_hdmi_in1_charsync0_ctl_pos_status[3:0];
assign vns_videooverlaysoc_csrbank6_data0_wer_value2_w = soc_videooverlaysoc_hdmi_in1_wer0_status[23:16];
assign vns_videooverlaysoc_csrbank6_data0_wer_value1_w = soc_videooverlaysoc_hdmi_in1_wer0_status[15:8];
assign vns_videooverlaysoc_csrbank6_data0_wer_value0_w = soc_videooverlaysoc_hdmi_in1_wer0_status[7:0];
assign vns_videooverlaysoc_csrbank6_data1_cap_phase_w = soc_videooverlaysoc_hdmi_in1_s7datacapture1_status[1:0];
assign vns_videooverlaysoc_csrbank6_data1_charsync_char_synced_w = soc_videooverlaysoc_hdmi_in1_charsync1_char_synced_status;
assign vns_videooverlaysoc_csrbank6_data1_charsync_ctl_pos_w = soc_videooverlaysoc_hdmi_in1_charsync1_ctl_pos_status[3:0];
assign vns_videooverlaysoc_csrbank6_data1_wer_value2_w = soc_videooverlaysoc_hdmi_in1_wer1_status[23:16];
assign vns_videooverlaysoc_csrbank6_data1_wer_value1_w = soc_videooverlaysoc_hdmi_in1_wer1_status[15:8];
assign vns_videooverlaysoc_csrbank6_data1_wer_value0_w = soc_videooverlaysoc_hdmi_in1_wer1_status[7:0];
assign vns_videooverlaysoc_csrbank6_data2_cap_phase_w = soc_videooverlaysoc_hdmi_in1_s7datacapture2_status[1:0];
assign vns_videooverlaysoc_csrbank6_data2_charsync_char_synced_w = soc_videooverlaysoc_hdmi_in1_charsync2_char_synced_status;
assign vns_videooverlaysoc_csrbank6_data2_charsync_ctl_pos_w = soc_videooverlaysoc_hdmi_in1_charsync2_ctl_pos_status[3:0];
assign vns_videooverlaysoc_csrbank6_data2_wer_value2_w = soc_videooverlaysoc_hdmi_in1_wer2_status[23:16];
assign vns_videooverlaysoc_csrbank6_data2_wer_value1_w = soc_videooverlaysoc_hdmi_in1_wer2_status[15:8];
assign vns_videooverlaysoc_csrbank6_data2_wer_value0_w = soc_videooverlaysoc_hdmi_in1_wer2_status[7:0];
assign vns_videooverlaysoc_csrbank6_chansync_channels_synced_w = soc_videooverlaysoc_hdmi_in1_chansync_status;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_storage = soc_videooverlaysoc_hdmi_in1_decode_terc4_storage_full;
assign vns_videooverlaysoc_csrbank6_decode_terc4_dvimode0_w = soc_videooverlaysoc_hdmi_in1_decode_terc4_storage_full;
assign vns_videooverlaysoc_csrbank6_resdetection_hres1_w = soc_videooverlaysoc_hdmi_in1_resdetection_hres_status[10:8];
assign vns_videooverlaysoc_csrbank6_resdetection_hres0_w = soc_videooverlaysoc_hdmi_in1_resdetection_hres_status[7:0];
assign vns_videooverlaysoc_csrbank6_resdetection_vres1_w = soc_videooverlaysoc_hdmi_in1_resdetection_vres_status[10:8];
assign vns_videooverlaysoc_csrbank6_resdetection_vres0_w = soc_videooverlaysoc_hdmi_in1_resdetection_vres_status[7:0];
assign soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage = soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full[28:5];
assign vns_videooverlaysoc_csrbank6_dma_frame_size3_w = soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full[28:24];
assign vns_videooverlaysoc_csrbank6_dma_frame_size2_w = soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full[23:16];
assign vns_videooverlaysoc_csrbank6_dma_frame_size1_w = soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full[15:8];
assign vns_videooverlaysoc_csrbank6_dma_frame_size0_w = {soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full[7:5], {3{1'd0}}};
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_storage = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_storage_full[1:0];
assign vns_videooverlaysoc_csrbank6_dma_slot0_status0_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_storage_full[1:0];
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[28:5];
assign vns_videooverlaysoc_csrbank6_dma_slot0_address3_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[28:24];
assign vns_videooverlaysoc_csrbank6_dma_slot0_address2_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[23:16];
assign vns_videooverlaysoc_csrbank6_dma_slot0_address1_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[15:8];
assign vns_videooverlaysoc_csrbank6_dma_slot0_address0_w = {soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[7:5], {3{1'd0}}};
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_storage = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_storage_full[1:0];
assign vns_videooverlaysoc_csrbank6_dma_slot1_status0_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_storage_full[1:0];
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[28:5];
assign vns_videooverlaysoc_csrbank6_dma_slot1_address3_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[28:24];
assign vns_videooverlaysoc_csrbank6_dma_slot1_address2_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[23:16];
assign vns_videooverlaysoc_csrbank6_dma_slot1_address1_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[15:8];
assign vns_videooverlaysoc_csrbank6_dma_slot1_address0_w = {soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[7:5], {3{1'd0}}};
assign soc_videooverlaysoc_hdmi_in1_dma_slot_array_storage = soc_videooverlaysoc_hdmi_in1_dma_slot_array_storage_full[1:0];
assign vns_videooverlaysoc_csrbank6_dma_ev_enable0_w = soc_videooverlaysoc_hdmi_in1_dma_slot_array_storage_full[1:0];
assign vns_videooverlaysoc_csrbank7_sel = (vns_videooverlaysoc_interface7_bank_bus_adr[13:9] == 5'd18);
assign vns_videooverlaysoc_csrbank7_value3_r = vns_videooverlaysoc_interface7_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank7_value3_re = ((vns_videooverlaysoc_csrbank7_sel & vns_videooverlaysoc_interface7_bank_bus_we) & (vns_videooverlaysoc_interface7_bank_bus_adr[1:0] == 1'd0));
assign vns_videooverlaysoc_csrbank7_value2_r = vns_videooverlaysoc_interface7_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank7_value2_re = ((vns_videooverlaysoc_csrbank7_sel & vns_videooverlaysoc_interface7_bank_bus_we) & (vns_videooverlaysoc_interface7_bank_bus_adr[1:0] == 1'd1));
assign vns_videooverlaysoc_csrbank7_value1_r = vns_videooverlaysoc_interface7_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank7_value1_re = ((vns_videooverlaysoc_csrbank7_sel & vns_videooverlaysoc_interface7_bank_bus_we) & (vns_videooverlaysoc_interface7_bank_bus_adr[1:0] == 2'd2));
assign vns_videooverlaysoc_csrbank7_value0_r = vns_videooverlaysoc_interface7_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank7_value0_re = ((vns_videooverlaysoc_csrbank7_sel & vns_videooverlaysoc_interface7_bank_bus_we) & (vns_videooverlaysoc_interface7_bank_bus_adr[1:0] == 2'd3));
assign vns_videooverlaysoc_csrbank7_value3_w = soc_videooverlaysoc_hdmi_in1_freq_status[31:24];
assign vns_videooverlaysoc_csrbank7_value2_w = soc_videooverlaysoc_hdmi_in1_freq_status[23:16];
assign vns_videooverlaysoc_csrbank7_value1_w = soc_videooverlaysoc_hdmi_in1_freq_status[15:8];
assign vns_videooverlaysoc_csrbank7_value0_w = soc_videooverlaysoc_hdmi_in1_freq_status[7:0];
assign vns_videooverlaysoc_csrbank8_sel = (vns_videooverlaysoc_interface8_bank_bus_adr[13:9] == 5'd22);
assign vns_videooverlaysoc_csrbank8_edid_snoop_adr0_r = vns_videooverlaysoc_interface8_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank8_edid_snoop_adr0_re = ((vns_videooverlaysoc_csrbank8_sel & vns_videooverlaysoc_interface8_bank_bus_we) & (vns_videooverlaysoc_interface8_bank_bus_adr[0] == 1'd0));
assign vns_videooverlaysoc_csrbank8_edid_snoop_dat_r = vns_videooverlaysoc_interface8_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank8_edid_snoop_dat_re = ((vns_videooverlaysoc_csrbank8_sel & vns_videooverlaysoc_interface8_bank_bus_we) & (vns_videooverlaysoc_interface8_bank_bus_adr[0] == 1'd1));
assign soc_videooverlaysoc_i2c_snoop_storage = soc_videooverlaysoc_i2c_snoop_storage_full[7:0];
assign vns_videooverlaysoc_csrbank8_edid_snoop_adr0_w = soc_videooverlaysoc_i2c_snoop_storage_full[7:0];
assign vns_videooverlaysoc_csrbank8_edid_snoop_dat_w = soc_videooverlaysoc_i2c_snoop_status[7:0];
assign vns_videooverlaysoc_sram2_sel = (vns_videooverlaysoc_interface2_sram_bus_adr[13:9] == 3'd4);
always @(*) begin
	vns_videooverlaysoc_interface2_sram_bus_dat_r <= 8'd0;
	if (vns_videooverlaysoc_sram2_sel_r) begin
		vns_videooverlaysoc_interface2_sram_bus_dat_r <= vns_videooverlaysoc_sram2_dat_r;
	end
end
assign vns_videooverlaysoc_sram2_adr = vns_videooverlaysoc_interface2_sram_bus_adr[4:0];
assign vns_videooverlaysoc_csrbank9_sel = (vns_videooverlaysoc_interface9_bank_bus_adr[13:9] == 5'd20);
assign vns_videooverlaysoc_csrbank9_hrect_start1_r = vns_videooverlaysoc_interface9_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank9_hrect_start1_re = ((vns_videooverlaysoc_csrbank9_sel & vns_videooverlaysoc_interface9_bank_bus_we) & (vns_videooverlaysoc_interface9_bank_bus_adr[3:0] == 1'd0));
assign vns_videooverlaysoc_csrbank9_hrect_start0_r = vns_videooverlaysoc_interface9_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank9_hrect_start0_re = ((vns_videooverlaysoc_csrbank9_sel & vns_videooverlaysoc_interface9_bank_bus_we) & (vns_videooverlaysoc_interface9_bank_bus_adr[3:0] == 1'd1));
assign vns_videooverlaysoc_csrbank9_hrect_end1_r = vns_videooverlaysoc_interface9_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank9_hrect_end1_re = ((vns_videooverlaysoc_csrbank9_sel & vns_videooverlaysoc_interface9_bank_bus_we) & (vns_videooverlaysoc_interface9_bank_bus_adr[3:0] == 2'd2));
assign vns_videooverlaysoc_csrbank9_hrect_end0_r = vns_videooverlaysoc_interface9_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank9_hrect_end0_re = ((vns_videooverlaysoc_csrbank9_sel & vns_videooverlaysoc_interface9_bank_bus_we) & (vns_videooverlaysoc_interface9_bank_bus_adr[3:0] == 2'd3));
assign vns_videooverlaysoc_csrbank9_vrect_start1_r = vns_videooverlaysoc_interface9_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank9_vrect_start1_re = ((vns_videooverlaysoc_csrbank9_sel & vns_videooverlaysoc_interface9_bank_bus_we) & (vns_videooverlaysoc_interface9_bank_bus_adr[3:0] == 3'd4));
assign vns_videooverlaysoc_csrbank9_vrect_start0_r = vns_videooverlaysoc_interface9_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank9_vrect_start0_re = ((vns_videooverlaysoc_csrbank9_sel & vns_videooverlaysoc_interface9_bank_bus_we) & (vns_videooverlaysoc_interface9_bank_bus_adr[3:0] == 3'd5));
assign vns_videooverlaysoc_csrbank9_vrect_end1_r = vns_videooverlaysoc_interface9_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank9_vrect_end1_re = ((vns_videooverlaysoc_csrbank9_sel & vns_videooverlaysoc_interface9_bank_bus_we) & (vns_videooverlaysoc_interface9_bank_bus_adr[3:0] == 3'd6));
assign vns_videooverlaysoc_csrbank9_vrect_end0_r = vns_videooverlaysoc_interface9_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank9_vrect_end0_re = ((vns_videooverlaysoc_csrbank9_sel & vns_videooverlaysoc_interface9_bank_bus_we) & (vns_videooverlaysoc_interface9_bank_bus_adr[3:0] == 3'd7));
assign vns_videooverlaysoc_csrbank9_rect_thresh0_r = vns_videooverlaysoc_interface9_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank9_rect_thresh0_re = ((vns_videooverlaysoc_csrbank9_sel & vns_videooverlaysoc_interface9_bank_bus_we) & (vns_videooverlaysoc_interface9_bank_bus_adr[3:0] == 4'd8));
assign soc_videooverlaysoc_hrect_start_storage = soc_videooverlaysoc_hrect_start_storage_full[11:0];
assign vns_videooverlaysoc_csrbank9_hrect_start1_w = soc_videooverlaysoc_hrect_start_storage_full[11:8];
assign vns_videooverlaysoc_csrbank9_hrect_start0_w = soc_videooverlaysoc_hrect_start_storage_full[7:0];
assign soc_videooverlaysoc_hrect_end_storage = soc_videooverlaysoc_hrect_end_storage_full[11:0];
assign vns_videooverlaysoc_csrbank9_hrect_end1_w = soc_videooverlaysoc_hrect_end_storage_full[11:8];
assign vns_videooverlaysoc_csrbank9_hrect_end0_w = soc_videooverlaysoc_hrect_end_storage_full[7:0];
assign soc_videooverlaysoc_vrect_start_storage = soc_videooverlaysoc_vrect_start_storage_full[11:0];
assign vns_videooverlaysoc_csrbank9_vrect_start1_w = soc_videooverlaysoc_vrect_start_storage_full[11:8];
assign vns_videooverlaysoc_csrbank9_vrect_start0_w = soc_videooverlaysoc_vrect_start_storage_full[7:0];
assign soc_videooverlaysoc_vrect_end_storage = soc_videooverlaysoc_vrect_end_storage_full[11:0];
assign vns_videooverlaysoc_csrbank9_vrect_end1_w = soc_videooverlaysoc_vrect_end_storage_full[11:8];
assign vns_videooverlaysoc_csrbank9_vrect_end0_w = soc_videooverlaysoc_vrect_end_storage_full[7:0];
assign soc_videooverlaysoc_rect_thresh_storage = soc_videooverlaysoc_rect_thresh_storage_full[7:0];
assign vns_videooverlaysoc_csrbank9_rect_thresh0_w = soc_videooverlaysoc_rect_thresh_storage_full[7:0];
assign vns_videooverlaysoc_csrbank10_sel = (vns_videooverlaysoc_interface10_bank_bus_adr[13:9] == 4'd8);
assign vns_videooverlaysoc_csrbank10_dfii_control0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank10_dfii_control0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 1'd0));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_command0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_command0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 1'd1));
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_issue_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_issue_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 2'd2));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_address1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_address1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 2'd3));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_address0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_address0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 3'd4));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_baddress0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[2:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_baddress0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 3'd5));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata7_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata7_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 3'd6));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata6_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata6_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 3'd7));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata5_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata5_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 4'd8));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata4_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata4_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 4'd9));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata3_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata3_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 4'd10));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata2_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata2_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 4'd11));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 4'd12));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 4'd13));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata7_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata7_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 4'd14));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata6_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata6_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 4'd15));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata5_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata5_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd16));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata4_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata4_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd17));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata3_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata3_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd18));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata2_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata2_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd19));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd20));
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd21));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_command0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_command0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd22));
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_issue_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_issue_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd23));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_address1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_address1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd24));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_address0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_address0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd25));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_baddress0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[2:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_baddress0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd26));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata7_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata7_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd27));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata6_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata6_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd28));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata5_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata5_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd29));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata4_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata4_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd30));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata3_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata3_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 5'd31));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata2_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata2_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd32));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd33));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd34));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata7_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata7_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd35));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata6_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata6_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd36));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata5_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata5_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd37));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata4_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata4_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd38));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata3_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata3_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd39));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata2_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata2_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd40));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd41));
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd42));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_command0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_command0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd43));
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_issue_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_issue_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd44));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_address1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_address1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd45));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_address0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_address0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd46));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_baddress0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[2:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_baddress0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd47));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata7_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata7_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd48));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata6_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata6_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd49));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata5_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata5_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd50));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata4_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata4_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd51));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata3_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata3_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd52));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata2_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata2_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd53));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd54));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd55));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata7_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata7_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd56));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata6_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata6_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd57));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata5_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata5_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd58));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata4_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata4_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd59));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata3_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata3_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd60));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata2_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata2_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd61));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd62));
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 6'd63));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_command0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_command0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd64));
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_issue_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_issue_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd65));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_address1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_address1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd66));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_address0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_address0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd67));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_baddress0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[2:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_baddress0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd68));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata7_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata7_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd69));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata6_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata6_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd70));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata5_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata5_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd71));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata4_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata4_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd72));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata3_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata3_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd73));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata2_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata2_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd74));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd75));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd76));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata7_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata7_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd77));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata6_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata6_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd78));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata5_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata5_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd79));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata4_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata4_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd80));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata3_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata3_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd81));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata2_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata2_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd82));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd83));
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd84));
assign soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_update_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_update_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd85));
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads2_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads2_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd86));
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd87));
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd88));
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites2_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites2_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd89));
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd90));
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd91));
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width1_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width1_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd92));
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width0_r = vns_videooverlaysoc_interface10_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width0_re = ((vns_videooverlaysoc_csrbank10_sel & vns_videooverlaysoc_interface10_bank_bus_we) & (vns_videooverlaysoc_interface10_bank_bus_adr[6:0] == 7'd93));
assign soc_videooverlaysoc_videooverlaysoc_sdram_storage = soc_videooverlaysoc_videooverlaysoc_sdram_storage_full[3:0];
assign vns_videooverlaysoc_csrbank10_dfii_control0_w = soc_videooverlaysoc_videooverlaysoc_sdram_storage_full[3:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage_full[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_command0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage_full[5:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_storage_full[13:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_address1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_storage_full[13:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_address0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_storage_full[7:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_storage_full[2:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_baddress0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_storage_full[2:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[63:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata7_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[63:56];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata6_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[55:48];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata5_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[47:40];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata4_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[39:32];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata3_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[31:24];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata2_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[23:16];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[15:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata7_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status[63:56];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata6_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status[55:48];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata5_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status[47:40];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata4_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status[39:32];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata3_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status[31:24];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata2_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status[23:16];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status[15:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi0_rddata0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status[7:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage_full[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_command0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage_full[5:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_storage_full[13:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_address1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_storage_full[13:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_address0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_storage_full[7:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_storage_full[2:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_baddress0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_storage_full[2:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[63:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata7_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[63:56];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata6_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[55:48];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata5_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[47:40];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata4_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[39:32];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata3_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[31:24];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata2_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[23:16];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[15:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata7_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status[63:56];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata6_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status[55:48];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata5_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status[47:40];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata4_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status[39:32];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata3_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status[31:24];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata2_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status[23:16];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status[15:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi1_rddata0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status[7:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage_full[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_command0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage_full[5:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_storage_full[13:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_address1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_storage_full[13:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_address0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_storage_full[7:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_storage_full[2:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_baddress0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_storage_full[2:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[63:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata7_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[63:56];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata6_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[55:48];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata5_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[47:40];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata4_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[39:32];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata3_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[31:24];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata2_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[23:16];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[15:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata7_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status[63:56];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata6_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status[55:48];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata5_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status[47:40];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata4_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status[39:32];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata3_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status[31:24];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata2_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status[23:16];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status[15:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi2_rddata0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status[7:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage_full[5:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_command0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage_full[5:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_storage_full[13:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_address1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_storage_full[13:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_address0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_storage_full[7:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_storage_full[2:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_baddress0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_storage_full[2:0];
assign soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[63:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata7_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[63:56];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata6_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[55:48];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata5_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[47:40];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata4_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[39:32];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata3_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[31:24];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata2_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[23:16];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[15:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[7:0];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata7_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status[63:56];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata6_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status[55:48];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata5_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status[47:40];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata4_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status[39:32];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata3_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status[31:24];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata2_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status[23:16];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata1_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status[15:8];
assign vns_videooverlaysoc_csrbank10_dfii_pi3_rddata0_w = soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status[7:0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads2_w = soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads_status[23:16];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads1_w = soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads_status[15:8];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads0_w = soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads_status[7:0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites2_w = soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites_status[23:16];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites1_w = soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites_status[15:8];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites0_w = soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites_status[7:0];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width1_w = soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_data_width_status[8];
assign vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width0_w = soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_data_width_status[7:0];
assign vns_videooverlaysoc_csrbank11_sel = (vns_videooverlaysoc_interface11_bank_bus_adr[13:9] == 3'd5);
assign vns_videooverlaysoc_csrbank11_load3_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_load3_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 1'd0));
assign vns_videooverlaysoc_csrbank11_load2_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_load2_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 1'd1));
assign vns_videooverlaysoc_csrbank11_load1_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_load1_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 2'd2));
assign vns_videooverlaysoc_csrbank11_load0_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_load0_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 2'd3));
assign vns_videooverlaysoc_csrbank11_reload3_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_reload3_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 3'd4));
assign vns_videooverlaysoc_csrbank11_reload2_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_reload2_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 3'd5));
assign vns_videooverlaysoc_csrbank11_reload1_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_reload1_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 3'd6));
assign vns_videooverlaysoc_csrbank11_reload0_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_reload0_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 3'd7));
assign vns_videooverlaysoc_csrbank11_en0_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank11_en0_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 4'd8));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_update_value_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_update_value_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 4'd9));
assign vns_videooverlaysoc_csrbank11_value3_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_value3_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 4'd10));
assign vns_videooverlaysoc_csrbank11_value2_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_value2_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 4'd11));
assign vns_videooverlaysoc_csrbank11_value1_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_value1_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 4'd12));
assign vns_videooverlaysoc_csrbank11_value0_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank11_value0_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 4'd13));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_status_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_status_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 4'd14));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_pending_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_pending_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 4'd15));
assign vns_videooverlaysoc_csrbank11_ev_enable0_r = vns_videooverlaysoc_interface11_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank11_ev_enable0_re = ((vns_videooverlaysoc_csrbank11_sel & vns_videooverlaysoc_interface11_bank_bus_we) & (vns_videooverlaysoc_interface11_bank_bus_adr[4:0] == 5'd16));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full[31:0];
assign vns_videooverlaysoc_csrbank11_load3_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full[31:24];
assign vns_videooverlaysoc_csrbank11_load2_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full[23:16];
assign vns_videooverlaysoc_csrbank11_load1_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full[15:8];
assign vns_videooverlaysoc_csrbank11_load0_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full[7:0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full[31:0];
assign vns_videooverlaysoc_csrbank11_reload3_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full[31:24];
assign vns_videooverlaysoc_csrbank11_reload2_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full[23:16];
assign vns_videooverlaysoc_csrbank11_reload1_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full[15:8];
assign vns_videooverlaysoc_csrbank11_reload0_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full[7:0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_storage = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_storage_full;
assign vns_videooverlaysoc_csrbank11_en0_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_storage_full;
assign vns_videooverlaysoc_csrbank11_value3_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value_status[31:24];
assign vns_videooverlaysoc_csrbank11_value2_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value_status[23:16];
assign vns_videooverlaysoc_csrbank11_value1_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value_status[15:8];
assign vns_videooverlaysoc_csrbank11_value0_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value_status[7:0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_storage = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_storage_full;
assign vns_videooverlaysoc_csrbank11_ev_enable0_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_storage_full;
assign vns_videooverlaysoc_csrbank12_sel = (vns_videooverlaysoc_interface12_bank_bus_adr[13:9] == 2'd3);
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxtx_r = vns_videooverlaysoc_interface12_bank_bus_dat_w[7:0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxtx_re = ((vns_videooverlaysoc_csrbank12_sel & vns_videooverlaysoc_interface12_bank_bus_we) & (vns_videooverlaysoc_interface12_bank_bus_adr[2:0] == 1'd0));
assign vns_videooverlaysoc_csrbank12_txfull_r = vns_videooverlaysoc_interface12_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank12_txfull_re = ((vns_videooverlaysoc_csrbank12_sel & vns_videooverlaysoc_interface12_bank_bus_we) & (vns_videooverlaysoc_interface12_bank_bus_adr[2:0] == 1'd1));
assign vns_videooverlaysoc_csrbank12_rxempty_r = vns_videooverlaysoc_interface12_bank_bus_dat_w[0];
assign vns_videooverlaysoc_csrbank12_rxempty_re = ((vns_videooverlaysoc_csrbank12_sel & vns_videooverlaysoc_interface12_bank_bus_we) & (vns_videooverlaysoc_interface12_bank_bus_adr[2:0] == 2'd2));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_status_r = vns_videooverlaysoc_interface12_bank_bus_dat_w[1:0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_status_re = ((vns_videooverlaysoc_csrbank12_sel & vns_videooverlaysoc_interface12_bank_bus_we) & (vns_videooverlaysoc_interface12_bank_bus_adr[2:0] == 2'd3));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_r = vns_videooverlaysoc_interface12_bank_bus_dat_w[1:0];
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_re = ((vns_videooverlaysoc_csrbank12_sel & vns_videooverlaysoc_interface12_bank_bus_we) & (vns_videooverlaysoc_interface12_bank_bus_adr[2:0] == 3'd4));
assign vns_videooverlaysoc_csrbank12_ev_enable0_r = vns_videooverlaysoc_interface12_bank_bus_dat_w[1:0];
assign vns_videooverlaysoc_csrbank12_ev_enable0_re = ((vns_videooverlaysoc_csrbank12_sel & vns_videooverlaysoc_interface12_bank_bus_we) & (vns_videooverlaysoc_interface12_bank_bus_adr[2:0] == 3'd5));
assign vns_videooverlaysoc_csrbank12_txfull_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_txfull_status;
assign vns_videooverlaysoc_csrbank12_rxempty_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxempty_status;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_storage = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_storage_full[1:0];
assign vns_videooverlaysoc_csrbank12_ev_enable0_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_storage_full[1:0];
assign vns_videooverlaysoc_csrbank13_sel = (vns_videooverlaysoc_interface13_bank_bus_adr[13:9] == 2'd2);
assign vns_videooverlaysoc_csrbank13_tuning_word3_r = vns_videooverlaysoc_interface13_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank13_tuning_word3_re = ((vns_videooverlaysoc_csrbank13_sel & vns_videooverlaysoc_interface13_bank_bus_we) & (vns_videooverlaysoc_interface13_bank_bus_adr[1:0] == 1'd0));
assign vns_videooverlaysoc_csrbank13_tuning_word2_r = vns_videooverlaysoc_interface13_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank13_tuning_word2_re = ((vns_videooverlaysoc_csrbank13_sel & vns_videooverlaysoc_interface13_bank_bus_we) & (vns_videooverlaysoc_interface13_bank_bus_adr[1:0] == 1'd1));
assign vns_videooverlaysoc_csrbank13_tuning_word1_r = vns_videooverlaysoc_interface13_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank13_tuning_word1_re = ((vns_videooverlaysoc_csrbank13_sel & vns_videooverlaysoc_interface13_bank_bus_we) & (vns_videooverlaysoc_interface13_bank_bus_adr[1:0] == 2'd2));
assign vns_videooverlaysoc_csrbank13_tuning_word0_r = vns_videooverlaysoc_interface13_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank13_tuning_word0_re = ((vns_videooverlaysoc_csrbank13_sel & vns_videooverlaysoc_interface13_bank_bus_we) & (vns_videooverlaysoc_interface13_bank_bus_adr[1:0] == 2'd3));
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full[31:0];
assign vns_videooverlaysoc_csrbank13_tuning_word3_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full[31:24];
assign vns_videooverlaysoc_csrbank13_tuning_word2_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full[23:16];
assign vns_videooverlaysoc_csrbank13_tuning_word1_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full[15:8];
assign vns_videooverlaysoc_csrbank13_tuning_word0_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full[7:0];
assign vns_videooverlaysoc_csrbank14_sel = (vns_videooverlaysoc_interface14_bank_bus_adr[13:9] == 4'd11);
assign vns_videooverlaysoc_csrbank14_temperature1_r = vns_videooverlaysoc_interface14_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank14_temperature1_re = ((vns_videooverlaysoc_csrbank14_sel & vns_videooverlaysoc_interface14_bank_bus_we) & (vns_videooverlaysoc_interface14_bank_bus_adr[2:0] == 1'd0));
assign vns_videooverlaysoc_csrbank14_temperature0_r = vns_videooverlaysoc_interface14_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank14_temperature0_re = ((vns_videooverlaysoc_csrbank14_sel & vns_videooverlaysoc_interface14_bank_bus_we) & (vns_videooverlaysoc_interface14_bank_bus_adr[2:0] == 1'd1));
assign vns_videooverlaysoc_csrbank14_vccint1_r = vns_videooverlaysoc_interface14_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank14_vccint1_re = ((vns_videooverlaysoc_csrbank14_sel & vns_videooverlaysoc_interface14_bank_bus_we) & (vns_videooverlaysoc_interface14_bank_bus_adr[2:0] == 2'd2));
assign vns_videooverlaysoc_csrbank14_vccint0_r = vns_videooverlaysoc_interface14_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank14_vccint0_re = ((vns_videooverlaysoc_csrbank14_sel & vns_videooverlaysoc_interface14_bank_bus_we) & (vns_videooverlaysoc_interface14_bank_bus_adr[2:0] == 2'd3));
assign vns_videooverlaysoc_csrbank14_vccaux1_r = vns_videooverlaysoc_interface14_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank14_vccaux1_re = ((vns_videooverlaysoc_csrbank14_sel & vns_videooverlaysoc_interface14_bank_bus_we) & (vns_videooverlaysoc_interface14_bank_bus_adr[2:0] == 3'd4));
assign vns_videooverlaysoc_csrbank14_vccaux0_r = vns_videooverlaysoc_interface14_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank14_vccaux0_re = ((vns_videooverlaysoc_csrbank14_sel & vns_videooverlaysoc_interface14_bank_bus_we) & (vns_videooverlaysoc_interface14_bank_bus_adr[2:0] == 3'd5));
assign vns_videooverlaysoc_csrbank14_vccbram1_r = vns_videooverlaysoc_interface14_bank_bus_dat_w[3:0];
assign vns_videooverlaysoc_csrbank14_vccbram1_re = ((vns_videooverlaysoc_csrbank14_sel & vns_videooverlaysoc_interface14_bank_bus_we) & (vns_videooverlaysoc_interface14_bank_bus_adr[2:0] == 3'd6));
assign vns_videooverlaysoc_csrbank14_vccbram0_r = vns_videooverlaysoc_interface14_bank_bus_dat_w[7:0];
assign vns_videooverlaysoc_csrbank14_vccbram0_re = ((vns_videooverlaysoc_csrbank14_sel & vns_videooverlaysoc_interface14_bank_bus_we) & (vns_videooverlaysoc_interface14_bank_bus_adr[2:0] == 3'd7));
assign vns_videooverlaysoc_csrbank14_temperature1_w = soc_videooverlaysoc_videooverlaysoc_temperature_status[11:8];
assign vns_videooverlaysoc_csrbank14_temperature0_w = soc_videooverlaysoc_videooverlaysoc_temperature_status[7:0];
assign vns_videooverlaysoc_csrbank14_vccint1_w = soc_videooverlaysoc_videooverlaysoc_vccint_status[11:8];
assign vns_videooverlaysoc_csrbank14_vccint0_w = soc_videooverlaysoc_videooverlaysoc_vccint_status[7:0];
assign vns_videooverlaysoc_csrbank14_vccaux1_w = soc_videooverlaysoc_videooverlaysoc_vccaux_status[11:8];
assign vns_videooverlaysoc_csrbank14_vccaux0_w = soc_videooverlaysoc_videooverlaysoc_vccaux_status[7:0];
assign vns_videooverlaysoc_csrbank14_vccbram1_w = soc_videooverlaysoc_videooverlaysoc_vccbram_status[11:8];
assign vns_videooverlaysoc_csrbank14_vccbram0_w = soc_videooverlaysoc_videooverlaysoc_vccbram_status[7:0];
assign vns_videooverlaysoc_interface0_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface1_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface2_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface3_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface4_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface5_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface6_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface7_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface8_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface9_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface10_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface11_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface12_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface13_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface14_bank_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface0_sram_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface1_sram_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface2_sram_bus_adr = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr;
assign vns_videooverlaysoc_interface0_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface1_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface2_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface3_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface4_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface5_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface6_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface7_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface8_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface9_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface10_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface11_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface12_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface13_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface14_bank_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface0_sram_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface1_sram_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface2_sram_bus_we = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we;
assign vns_videooverlaysoc_interface0_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface1_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface2_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface3_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface4_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface5_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface6_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface7_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface8_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface9_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface10_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface11_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface12_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface13_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface14_bank_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface0_sram_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface1_sram_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign vns_videooverlaysoc_interface2_sram_bus_dat_w = soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_r = (((((((((((((((((vns_videooverlaysoc_interface0_bank_bus_dat_r | vns_videooverlaysoc_interface1_bank_bus_dat_r) | vns_videooverlaysoc_interface2_bank_bus_dat_r) | vns_videooverlaysoc_interface3_bank_bus_dat_r) | vns_videooverlaysoc_interface4_bank_bus_dat_r) | vns_videooverlaysoc_interface5_bank_bus_dat_r) | vns_videooverlaysoc_interface6_bank_bus_dat_r) | vns_videooverlaysoc_interface7_bank_bus_dat_r) | vns_videooverlaysoc_interface8_bank_bus_dat_r) | vns_videooverlaysoc_interface9_bank_bus_dat_r) | vns_videooverlaysoc_interface10_bank_bus_dat_r) | vns_videooverlaysoc_interface11_bank_bus_dat_r) | vns_videooverlaysoc_interface12_bank_bus_dat_r) | vns_videooverlaysoc_interface13_bank_bus_dat_r) | vns_videooverlaysoc_interface14_bank_bus_dat_r) | vns_videooverlaysoc_interface0_sram_bus_dat_r) | vns_videooverlaysoc_interface1_sram_bus_dat_r) | vns_videooverlaysoc_interface2_sram_bus_dat_r);
assign vns_slice_proxy0 = soc_videooverlaysoc_core_mac_depacketizer_header[111:96];
assign vns_slice_proxy1 = soc_videooverlaysoc_core_mac_depacketizer_header[111:96];
assign vns_slice_proxy2 = soc_videooverlaysoc_core_mac_depacketizer_header[95:48];
assign vns_slice_proxy3 = soc_videooverlaysoc_core_mac_depacketizer_header[95:48];
assign vns_slice_proxy4 = soc_videooverlaysoc_core_mac_depacketizer_header[95:48];
assign vns_slice_proxy5 = soc_videooverlaysoc_core_mac_depacketizer_header[95:48];
assign vns_slice_proxy6 = soc_videooverlaysoc_core_mac_depacketizer_header[95:48];
assign vns_slice_proxy7 = soc_videooverlaysoc_core_mac_depacketizer_header[95:48];
assign vns_slice_proxy8 = soc_videooverlaysoc_core_mac_depacketizer_header[47:0];
assign vns_slice_proxy9 = soc_videooverlaysoc_core_mac_depacketizer_header[47:0];
assign vns_slice_proxy10 = soc_videooverlaysoc_core_mac_depacketizer_header[47:0];
assign vns_slice_proxy11 = soc_videooverlaysoc_core_mac_depacketizer_header[47:0];
assign vns_slice_proxy12 = soc_videooverlaysoc_core_mac_depacketizer_header[47:0];
assign vns_slice_proxy13 = soc_videooverlaysoc_core_mac_depacketizer_header[47:0];
assign vns_slice_proxy14 = soc_videooverlaysoc_core_arp_depacketizer_header[39:32];
assign vns_slice_proxy15 = soc_videooverlaysoc_core_arp_depacketizer_header[15:0];
assign vns_slice_proxy16 = soc_videooverlaysoc_core_arp_depacketizer_header[15:0];
assign vns_slice_proxy17 = soc_videooverlaysoc_core_arp_depacketizer_header[63:48];
assign vns_slice_proxy18 = soc_videooverlaysoc_core_arp_depacketizer_header[63:48];
assign vns_slice_proxy19 = soc_videooverlaysoc_core_arp_depacketizer_header[31:16];
assign vns_slice_proxy20 = soc_videooverlaysoc_core_arp_depacketizer_header[31:16];
assign vns_slice_proxy21 = soc_videooverlaysoc_core_arp_depacketizer_header[47:40];
assign vns_slice_proxy22 = soc_videooverlaysoc_core_arp_depacketizer_header[143:112];
assign vns_slice_proxy23 = soc_videooverlaysoc_core_arp_depacketizer_header[143:112];
assign vns_slice_proxy24 = soc_videooverlaysoc_core_arp_depacketizer_header[143:112];
assign vns_slice_proxy25 = soc_videooverlaysoc_core_arp_depacketizer_header[143:112];
assign vns_slice_proxy26 = soc_videooverlaysoc_core_arp_depacketizer_header[111:64];
assign vns_slice_proxy27 = soc_videooverlaysoc_core_arp_depacketizer_header[111:64];
assign vns_slice_proxy28 = soc_videooverlaysoc_core_arp_depacketizer_header[111:64];
assign vns_slice_proxy29 = soc_videooverlaysoc_core_arp_depacketizer_header[111:64];
assign vns_slice_proxy30 = soc_videooverlaysoc_core_arp_depacketizer_header[111:64];
assign vns_slice_proxy31 = soc_videooverlaysoc_core_arp_depacketizer_header[111:64];
assign vns_slice_proxy32 = soc_videooverlaysoc_core_arp_depacketizer_header[223:192];
assign vns_slice_proxy33 = soc_videooverlaysoc_core_arp_depacketizer_header[223:192];
assign vns_slice_proxy34 = soc_videooverlaysoc_core_arp_depacketizer_header[223:192];
assign vns_slice_proxy35 = soc_videooverlaysoc_core_arp_depacketizer_header[223:192];
assign vns_slice_proxy36 = soc_videooverlaysoc_core_arp_depacketizer_header[191:144];
assign vns_slice_proxy37 = soc_videooverlaysoc_core_arp_depacketizer_header[191:144];
assign vns_slice_proxy38 = soc_videooverlaysoc_core_arp_depacketizer_header[191:144];
assign vns_slice_proxy39 = soc_videooverlaysoc_core_arp_depacketizer_header[191:144];
assign vns_slice_proxy40 = soc_videooverlaysoc_core_arp_depacketizer_header[191:144];
assign vns_slice_proxy41 = soc_videooverlaysoc_core_arp_depacketizer_header[191:144];
assign vns_slice_proxy42 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[95:80];
assign vns_slice_proxy43 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[95:80];
assign vns_slice_proxy44 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[47:32];
assign vns_slice_proxy45 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[47:32];
assign vns_slice_proxy46 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[3:0];
assign vns_slice_proxy47 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[79:72];
assign vns_slice_proxy48 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[127:96];
assign vns_slice_proxy49 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[127:96];
assign vns_slice_proxy50 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[127:96];
assign vns_slice_proxy51 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[127:96];
assign vns_slice_proxy52 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[159:128];
assign vns_slice_proxy53 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[159:128];
assign vns_slice_proxy54 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[159:128];
assign vns_slice_proxy55 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[159:128];
assign vns_slice_proxy56 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[31:16];
assign vns_slice_proxy57 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[31:16];
assign vns_slice_proxy58 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[71:64];
assign vns_slice_proxy59 = soc_videooverlaysoc_core_ip_rx_depacketizer_header[7:4];
assign vns_slice_proxy60 = soc_videooverlaysoc_core_icmp_rx_depacketizer_header[31:16];
assign vns_slice_proxy61 = soc_videooverlaysoc_core_icmp_rx_depacketizer_header[31:16];
assign vns_slice_proxy62 = soc_videooverlaysoc_core_icmp_rx_depacketizer_header[15:8];
assign vns_slice_proxy63 = soc_videooverlaysoc_core_icmp_rx_depacketizer_header[7:0];
assign vns_slice_proxy64 = soc_videooverlaysoc_core_icmp_rx_depacketizer_header[63:32];
assign vns_slice_proxy65 = soc_videooverlaysoc_core_icmp_rx_depacketizer_header[63:32];
assign vns_slice_proxy66 = soc_videooverlaysoc_core_icmp_rx_depacketizer_header[63:32];
assign vns_slice_proxy67 = soc_videooverlaysoc_core_icmp_rx_depacketizer_header[63:32];
assign vns_slice_proxy68 = soc_videooverlaysoc_core_depacketizer_header[63:48];
assign vns_slice_proxy69 = soc_videooverlaysoc_core_depacketizer_header[63:48];
assign vns_slice_proxy70 = soc_videooverlaysoc_core_depacketizer_header[31:16];
assign vns_slice_proxy71 = soc_videooverlaysoc_core_depacketizer_header[31:16];
assign vns_slice_proxy72 = soc_videooverlaysoc_core_depacketizer_header[47:32];
assign vns_slice_proxy73 = soc_videooverlaysoc_core_depacketizer_header[47:32];
assign vns_slice_proxy74 = soc_videooverlaysoc_core_depacketizer_header[15:0];
assign vns_slice_proxy75 = soc_videooverlaysoc_core_depacketizer_header[15:0];
assign vns_slice_proxy76 = soc_videooverlaysoc_packet_depacketizer_header[31:28];
assign vns_slice_proxy77 = soc_videooverlaysoc_packet_depacketizer_header[15:0];
assign vns_slice_proxy78 = soc_videooverlaysoc_packet_depacketizer_header[15:0];
assign vns_slice_proxy79 = soc_videooverlaysoc_packet_depacketizer_header[18];
assign vns_slice_proxy80 = soc_videooverlaysoc_packet_depacketizer_header[16];
assign vns_slice_proxy81 = soc_videooverlaysoc_packet_depacketizer_header[27:24];
assign vns_slice_proxy82 = soc_videooverlaysoc_packet_depacketizer_header[17];
assign vns_slice_proxy83 = soc_videooverlaysoc_packet_depacketizer_header[23:20];
assign vns_slice_proxy84 = soc_videooverlaysoc_record_depacketizer_header[0];
assign vns_slice_proxy85 = soc_videooverlaysoc_record_depacketizer_header[15:8];
assign vns_slice_proxy86 = soc_videooverlaysoc_record_depacketizer_header[4];
assign vns_slice_proxy87 = soc_videooverlaysoc_record_depacketizer_header[1];
assign vns_slice_proxy88 = soc_videooverlaysoc_record_depacketizer_header[31:24];
assign vns_slice_proxy89 = soc_videooverlaysoc_record_depacketizer_header[2];
assign vns_slice_proxy90 = soc_videooverlaysoc_record_depacketizer_header[5];
assign vns_slice_proxy91 = soc_videooverlaysoc_record_depacketizer_header[23:16];
assign vns_slice_proxy92 = soc_videooverlaysoc_record_depacketizer_header[6];
always @(*) begin
	vns_comb_rhs_array_muxed0 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[0];
		end
		1'd1: begin
			vns_comb_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[1];
		end
		2'd2: begin
			vns_comb_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[2];
		end
		2'd3: begin
			vns_comb_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[3];
		end
		3'd4: begin
			vns_comb_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[4];
		end
		3'd5: begin
			vns_comb_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[5];
		end
		3'd6: begin
			vns_comb_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[6];
		end
		default: begin
			vns_comb_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_valids[7];
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed1 <= 14'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_a;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_a;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_a;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_a;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_a;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_a;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_a;
		end
		default: begin
			vns_comb_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed2 <= 3'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ba;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ba;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ba;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ba;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ba;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ba;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ba;
		end
		default: begin
			vns_comb_rhs_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed3 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_read;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_read;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_read;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_read;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_read;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_read;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_read;
		end
		default: begin
			vns_comb_rhs_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_read;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed4 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_write;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_write;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_write;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_write;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_write;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_write;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_write;
		end
		default: begin
			vns_comb_rhs_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_write;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed5 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_cmd;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_cmd;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_cmd;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_cmd;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_cmd;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_cmd;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_cmd;
		end
		default: begin
			vns_comb_rhs_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_cmd;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed0 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_t_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_cas;
		end
		1'd1: begin
			vns_comb_t_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_cas;
		end
		2'd2: begin
			vns_comb_t_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_cas;
		end
		2'd3: begin
			vns_comb_t_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_cas;
		end
		3'd4: begin
			vns_comb_t_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_cas;
		end
		3'd5: begin
			vns_comb_t_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_cas;
		end
		3'd6: begin
			vns_comb_t_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_cas;
		end
		default: begin
			vns_comb_t_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed1 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_t_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ras;
		end
		1'd1: begin
			vns_comb_t_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ras;
		end
		2'd2: begin
			vns_comb_t_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ras;
		end
		2'd3: begin
			vns_comb_t_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ras;
		end
		3'd4: begin
			vns_comb_t_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ras;
		end
		3'd5: begin
			vns_comb_t_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ras;
		end
		3'd6: begin
			vns_comb_t_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ras;
		end
		default: begin
			vns_comb_t_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed2 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_t_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_t_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_we;
		end
		2'd2: begin
			vns_comb_t_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_we;
		end
		2'd3: begin
			vns_comb_t_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_we;
		end
		3'd4: begin
			vns_comb_t_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_we;
		end
		3'd5: begin
			vns_comb_t_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_we;
		end
		3'd6: begin
			vns_comb_t_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_we;
		end
		default: begin
			vns_comb_t_array_muxed2 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed6 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed6 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[0];
		end
		1'd1: begin
			vns_comb_rhs_array_muxed6 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[1];
		end
		2'd2: begin
			vns_comb_rhs_array_muxed6 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[2];
		end
		2'd3: begin
			vns_comb_rhs_array_muxed6 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[3];
		end
		3'd4: begin
			vns_comb_rhs_array_muxed6 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[4];
		end
		3'd5: begin
			vns_comb_rhs_array_muxed6 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[5];
		end
		3'd6: begin
			vns_comb_rhs_array_muxed6 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[6];
		end
		default: begin
			vns_comb_rhs_array_muxed6 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_valids[7];
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed7 <= 14'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_a;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_a;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_a;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_a;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_a;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_a;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_a;
		end
		default: begin
			vns_comb_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed8 <= 3'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ba;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ba;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ba;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ba;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ba;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ba;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ba;
		end
		default: begin
			vns_comb_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed9 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed9 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_read;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed9 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_read;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed9 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_read;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed9 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_read;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed9 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_read;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed9 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_read;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed9 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_read;
		end
		default: begin
			vns_comb_rhs_array_muxed9 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_read;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed10 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed10 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_write;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed10 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_write;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed10 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_write;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed10 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_write;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed10 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_write;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed10 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_write;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed10 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_write;
		end
		default: begin
			vns_comb_rhs_array_muxed10 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_write;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed11 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed11 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_is_cmd;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed11 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_is_cmd;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed11 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_is_cmd;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed11 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_is_cmd;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed11 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_is_cmd;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed11 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_is_cmd;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed11 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_is_cmd;
		end
		default: begin
			vns_comb_rhs_array_muxed11 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_is_cmd;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed3 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_t_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_cas;
		end
		1'd1: begin
			vns_comb_t_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_cas;
		end
		2'd2: begin
			vns_comb_t_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_cas;
		end
		2'd3: begin
			vns_comb_t_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_cas;
		end
		3'd4: begin
			vns_comb_t_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_cas;
		end
		3'd5: begin
			vns_comb_t_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_cas;
		end
		3'd6: begin
			vns_comb_t_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_cas;
		end
		default: begin
			vns_comb_t_array_muxed3 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed4 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_t_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_ras;
		end
		1'd1: begin
			vns_comb_t_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_ras;
		end
		2'd2: begin
			vns_comb_t_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_ras;
		end
		2'd3: begin
			vns_comb_t_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_ras;
		end
		3'd4: begin
			vns_comb_t_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_ras;
		end
		3'd5: begin
			vns_comb_t_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_ras;
		end
		3'd6: begin
			vns_comb_t_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_ras;
		end
		default: begin
			vns_comb_t_array_muxed4 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed5 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_t_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_t_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_payload_we;
		end
		2'd2: begin
			vns_comb_t_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_payload_we;
		end
		2'd3: begin
			vns_comb_t_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_payload_we;
		end
		3'd4: begin
			vns_comb_t_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_payload_we;
		end
		3'd5: begin
			vns_comb_t_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_payload_we;
		end
		3'd6: begin
			vns_comb_t_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_payload_we;
		end
		default: begin
			vns_comb_t_array_muxed5 <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed12 <= 21'd0;
	case (vns_roundrobin0_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed12 <= {soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[23:10], soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[6:0]};
		end
		1'd1: begin
			vns_comb_rhs_array_muxed12 <= {soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[23:10], soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[6:0]};
		end
		default: begin
			vns_comb_rhs_array_muxed12 <= {soc_videooverlaysoc_out_dram_port_cmd_payload_addr[23:10], soc_videooverlaysoc_out_dram_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed13 <= 1'd0;
	case (vns_roundrobin0_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed13 <= soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed13 <= soc_videooverlaysoc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed13 <= soc_videooverlaysoc_out_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed14 <= 1'd0;
	case (vns_roundrobin0_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed14 <= (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 1'd0) & (~(((((((vns_locked0 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed14 <= (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 1'd0) & (~(((((((vns_locked1 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed14 <= (((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 1'd0) & (~(((((((vns_locked2 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed15 <= 21'd0;
	case (vns_roundrobin1_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed15 <= {soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[23:10], soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[6:0]};
		end
		1'd1: begin
			vns_comb_rhs_array_muxed15 <= {soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[23:10], soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[6:0]};
		end
		default: begin
			vns_comb_rhs_array_muxed15 <= {soc_videooverlaysoc_out_dram_port_cmd_payload_addr[23:10], soc_videooverlaysoc_out_dram_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed16 <= 1'd0;
	case (vns_roundrobin1_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed16 <= soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed16 <= soc_videooverlaysoc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed16 <= soc_videooverlaysoc_out_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed17 <= 1'd0;
	case (vns_roundrobin1_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed17 <= (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 1'd1) & (~(((((((vns_locked3 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed17 <= (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 1'd1) & (~(((((((vns_locked4 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed17 <= (((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 1'd1) & (~(((((((vns_locked5 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed18 <= 21'd0;
	case (vns_roundrobin2_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed18 <= {soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[23:10], soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[6:0]};
		end
		1'd1: begin
			vns_comb_rhs_array_muxed18 <= {soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[23:10], soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[6:0]};
		end
		default: begin
			vns_comb_rhs_array_muxed18 <= {soc_videooverlaysoc_out_dram_port_cmd_payload_addr[23:10], soc_videooverlaysoc_out_dram_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed19 <= 1'd0;
	case (vns_roundrobin2_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed19 <= soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed19 <= soc_videooverlaysoc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed19 <= soc_videooverlaysoc_out_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed20 <= 1'd0;
	case (vns_roundrobin2_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed20 <= (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 2'd2) & (~(((((((vns_locked6 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed20 <= (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 2'd2) & (~(((((((vns_locked7 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed20 <= (((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 2'd2) & (~(((((((vns_locked8 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed21 <= 21'd0;
	case (vns_roundrobin3_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed21 <= {soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[23:10], soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[6:0]};
		end
		1'd1: begin
			vns_comb_rhs_array_muxed21 <= {soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[23:10], soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[6:0]};
		end
		default: begin
			vns_comb_rhs_array_muxed21 <= {soc_videooverlaysoc_out_dram_port_cmd_payload_addr[23:10], soc_videooverlaysoc_out_dram_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed22 <= 1'd0;
	case (vns_roundrobin3_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed22 <= soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed22 <= soc_videooverlaysoc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed22 <= soc_videooverlaysoc_out_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed23 <= 1'd0;
	case (vns_roundrobin3_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed23 <= (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 2'd3) & (~(((((((vns_locked9 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed23 <= (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 2'd3) & (~(((((((vns_locked10 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed23 <= (((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 2'd3) & (~(((((((vns_locked11 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed24 <= 21'd0;
	case (vns_roundrobin4_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed24 <= {soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[23:10], soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[6:0]};
		end
		1'd1: begin
			vns_comb_rhs_array_muxed24 <= {soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[23:10], soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[6:0]};
		end
		default: begin
			vns_comb_rhs_array_muxed24 <= {soc_videooverlaysoc_out_dram_port_cmd_payload_addr[23:10], soc_videooverlaysoc_out_dram_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed25 <= 1'd0;
	case (vns_roundrobin4_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed25 <= soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed25 <= soc_videooverlaysoc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed25 <= soc_videooverlaysoc_out_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed26 <= 1'd0;
	case (vns_roundrobin4_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed26 <= (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd4) & (~(((((((vns_locked12 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed26 <= (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd4) & (~(((((((vns_locked13 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed26 <= (((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd4) & (~(((((((vns_locked14 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed27 <= 21'd0;
	case (vns_roundrobin5_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed27 <= {soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[23:10], soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[6:0]};
		end
		1'd1: begin
			vns_comb_rhs_array_muxed27 <= {soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[23:10], soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[6:0]};
		end
		default: begin
			vns_comb_rhs_array_muxed27 <= {soc_videooverlaysoc_out_dram_port_cmd_payload_addr[23:10], soc_videooverlaysoc_out_dram_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed28 <= 1'd0;
	case (vns_roundrobin5_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed28 <= soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed28 <= soc_videooverlaysoc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed28 <= soc_videooverlaysoc_out_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed29 <= 1'd0;
	case (vns_roundrobin5_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed29 <= (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd5) & (~(((((((vns_locked15 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed29 <= (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd5) & (~(((((((vns_locked16 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed29 <= (((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd5) & (~(((((((vns_locked17 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed30 <= 21'd0;
	case (vns_roundrobin6_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed30 <= {soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[23:10], soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[6:0]};
		end
		1'd1: begin
			vns_comb_rhs_array_muxed30 <= {soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[23:10], soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[6:0]};
		end
		default: begin
			vns_comb_rhs_array_muxed30 <= {soc_videooverlaysoc_out_dram_port_cmd_payload_addr[23:10], soc_videooverlaysoc_out_dram_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed31 <= 1'd0;
	case (vns_roundrobin6_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed31 <= soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed31 <= soc_videooverlaysoc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed31 <= soc_videooverlaysoc_out_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed32 <= 1'd0;
	case (vns_roundrobin6_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed32 <= (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd6) & (~(((((((vns_locked18 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed32 <= (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd6) & (~(((((((vns_locked19 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed32 <= (((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd6) & (~(((((((vns_locked20 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed33 <= 21'd0;
	case (vns_roundrobin7_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed33 <= {soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[23:10], soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[6:0]};
		end
		1'd1: begin
			vns_comb_rhs_array_muxed33 <= {soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[23:10], soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[6:0]};
		end
		default: begin
			vns_comb_rhs_array_muxed33 <= {soc_videooverlaysoc_out_dram_port_cmd_payload_addr[23:10], soc_videooverlaysoc_out_dram_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed34 <= 1'd0;
	case (vns_roundrobin7_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed34 <= soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed34 <= soc_videooverlaysoc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed34 <= soc_videooverlaysoc_out_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed35 <= 1'd0;
	case (vns_roundrobin7_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed35 <= (((soc_videooverlaysoc_videooverlaysoc_port_cmd_payload_addr[9:7] == 3'd7) & (~(((((((vns_locked21 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))))) & soc_videooverlaysoc_videooverlaysoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed35 <= (((soc_videooverlaysoc_litedramcrossbar_cmd_payload_addr[9:7] == 3'd7) & (~(((((((vns_locked22 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))))) & soc_videooverlaysoc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed35 <= (((soc_videooverlaysoc_out_dram_port_cmd_payload_addr[9:7] == 3'd7) & (~(((((((vns_locked23 | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))))) & soc_videooverlaysoc_out_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed36 <= 24'd0;
	case (soc_videooverlaysoc_hdmi_in1_dma_slot_array_current_slot)
		1'd0: begin
			vns_comb_rhs_array_muxed36 <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address;
		end
		default: begin
			vns_comb_rhs_array_muxed36 <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed37 <= 1'd0;
	case (soc_videooverlaysoc_hdmi_in1_dma_slot_array_current_slot)
		1'd0: begin
			vns_comb_rhs_array_muxed37 <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_valid;
		end
		default: begin
			vns_comb_rhs_array_muxed37 <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_valid;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed38 <= 30'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed38 <= soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_adr;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed39 <= 32'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed39 <= soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_dat_w;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed40 <= 4'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed40 <= soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_sel;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed41 <= 1'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed41 <= soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_cyc;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed42 <= 1'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed42 <= soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_stb;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed43 <= 1'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed43 <= soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed44 <= 3'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed44 <= soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_cti;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed45 <= 2'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed45 <= soc_videooverlaysoc_videooverlaysoc_interface1_wb_sdram_bte;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed46 <= 30'd0;
	case (vns_videooverlaysoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed46 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_adr;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed46 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_adr;
		end
		default: begin
			vns_comb_rhs_array_muxed46 <= soc_videooverlaysoc_wishbone_bus_adr;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed47 <= 32'd0;
	case (vns_videooverlaysoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed47 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_dat_w;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed47 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_dat_w;
		end
		default: begin
			vns_comb_rhs_array_muxed47 <= soc_videooverlaysoc_wishbone_bus_dat_w;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed48 <= 4'd0;
	case (vns_videooverlaysoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed48 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_sel;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed48 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_sel;
		end
		default: begin
			vns_comb_rhs_array_muxed48 <= soc_videooverlaysoc_wishbone_bus_sel;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed49 <= 1'd0;
	case (vns_videooverlaysoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed49 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_cyc;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed49 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_cyc;
		end
		default: begin
			vns_comb_rhs_array_muxed49 <= soc_videooverlaysoc_wishbone_bus_cyc;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed50 <= 1'd0;
	case (vns_videooverlaysoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed50 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_stb;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed50 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_stb;
		end
		default: begin
			vns_comb_rhs_array_muxed50 <= soc_videooverlaysoc_wishbone_bus_stb;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed51 <= 1'd0;
	case (vns_videooverlaysoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed51 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed51 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_we;
		end
		default: begin
			vns_comb_rhs_array_muxed51 <= soc_videooverlaysoc_wishbone_bus_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed52 <= 3'd0;
	case (vns_videooverlaysoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed52 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_cti;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed52 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_cti;
		end
		default: begin
			vns_comb_rhs_array_muxed52 <= soc_videooverlaysoc_wishbone_bus_cti;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed53 <= 2'd0;
	case (vns_videooverlaysoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed53 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_bte;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed53 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_bte;
		end
		default: begin
			vns_comb_rhs_array_muxed53 <= soc_videooverlaysoc_wishbone_bus_bte;
		end
	endcase
end
always @(*) begin
	vns_sync_f_array_muxed0 <= 10'd0;
	case (soc_videooverlaysoc_encoder0_new_c2)
		1'd0: begin
			vns_sync_f_array_muxed0 <= 10'd852;
		end
		1'd1: begin
			vns_sync_f_array_muxed0 <= 8'd171;
		end
		2'd2: begin
			vns_sync_f_array_muxed0 <= 9'd340;
		end
		default: begin
			vns_sync_f_array_muxed0 <= 10'd683;
		end
	endcase
end
always @(*) begin
	vns_sync_f_array_muxed1 <= 10'd0;
	case (soc_videooverlaysoc_encoder1_new_c2)
		1'd0: begin
			vns_sync_f_array_muxed1 <= 10'd852;
		end
		1'd1: begin
			vns_sync_f_array_muxed1 <= 8'd171;
		end
		2'd2: begin
			vns_sync_f_array_muxed1 <= 9'd340;
		end
		default: begin
			vns_sync_f_array_muxed1 <= 10'd683;
		end
	endcase
end
always @(*) begin
	vns_sync_f_array_muxed2 <= 10'd0;
	case (soc_videooverlaysoc_encoder2_new_c2)
		1'd0: begin
			vns_sync_f_array_muxed2 <= 10'd852;
		end
		1'd1: begin
			vns_sync_f_array_muxed2 <= 8'd171;
		end
		2'd2: begin
			vns_sync_f_array_muxed2 <= 9'd340;
		end
		default: begin
			vns_sync_f_array_muxed2 <= 10'd683;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed0 <= 3'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_nop_ba[2:0];
		end
		1'd1: begin
			vns_sync_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ba[2:0];
		end
		2'd2: begin
			vns_sync_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ba[2:0];
		end
		default: begin
			vns_sync_rhs_array_muxed0 <= soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ba[2:0];
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed1 <= 14'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_nop_a;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			vns_sync_rhs_array_muxed1 <= soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed2 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed2 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed2 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed2 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_cas);
		end
		default: begin
			vns_sync_rhs_array_muxed2 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_cas);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed3 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed3 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed3 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed3 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ras);
		end
		default: begin
			vns_sync_rhs_array_muxed3 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ras);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed4 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed4 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed4 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed4 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_we);
		end
		default: begin
			vns_sync_rhs_array_muxed4 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_we);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed5 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed5 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed5 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed5 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			vns_sync_rhs_array_muxed5 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed6 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed6 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed6 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed6 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			vns_sync_rhs_array_muxed6 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed7 <= 3'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_nop_ba[2:0];
		end
		1'd1: begin
			vns_sync_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ba[2:0];
		end
		2'd2: begin
			vns_sync_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ba[2:0];
		end
		default: begin
			vns_sync_rhs_array_muxed7 <= soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ba[2:0];
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed8 <= 14'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_nop_a;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			vns_sync_rhs_array_muxed8 <= soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed9 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed9 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed9 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed9 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_cas);
		end
		default: begin
			vns_sync_rhs_array_muxed9 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_cas);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed10 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed10 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed10 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed10 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ras);
		end
		default: begin
			vns_sync_rhs_array_muxed10 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ras);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed11 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed11 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed11 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed11 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_we);
		end
		default: begin
			vns_sync_rhs_array_muxed11 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_we);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed12 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed12 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed12 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed12 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			vns_sync_rhs_array_muxed12 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed13 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed13 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed13 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed13 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			vns_sync_rhs_array_muxed13 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed14 <= 3'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed14 <= soc_videooverlaysoc_videooverlaysoc_sdram_nop_ba[2:0];
		end
		1'd1: begin
			vns_sync_rhs_array_muxed14 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ba[2:0];
		end
		2'd2: begin
			vns_sync_rhs_array_muxed14 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ba[2:0];
		end
		default: begin
			vns_sync_rhs_array_muxed14 <= soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ba[2:0];
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed15 <= 14'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed15 <= soc_videooverlaysoc_videooverlaysoc_sdram_nop_a;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed15 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed15 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			vns_sync_rhs_array_muxed15 <= soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed16 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed16 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed16 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed16 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_cas);
		end
		default: begin
			vns_sync_rhs_array_muxed16 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_cas);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed17 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed17 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed17 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed17 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ras);
		end
		default: begin
			vns_sync_rhs_array_muxed17 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ras);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed18 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed18 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed18 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed18 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_we);
		end
		default: begin
			vns_sync_rhs_array_muxed18 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_we);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed19 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed19 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed19 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed19 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			vns_sync_rhs_array_muxed19 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed20 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed20 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed20 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed20 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			vns_sync_rhs_array_muxed20 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed21 <= 3'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed21 <= soc_videooverlaysoc_videooverlaysoc_sdram_nop_ba[2:0];
		end
		1'd1: begin
			vns_sync_rhs_array_muxed21 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ba[2:0];
		end
		2'd2: begin
			vns_sync_rhs_array_muxed21 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ba[2:0];
		end
		default: begin
			vns_sync_rhs_array_muxed21 <= soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ba[2:0];
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed22 <= 14'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed22 <= soc_videooverlaysoc_videooverlaysoc_sdram_nop_a;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed22 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed22 <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			vns_sync_rhs_array_muxed22 <= soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed23 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed23 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed23 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_cas);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed23 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_cas);
		end
		default: begin
			vns_sync_rhs_array_muxed23 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_cas);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed24 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed24 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed24 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_ras);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed24 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_ras);
		end
		default: begin
			vns_sync_rhs_array_muxed24 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ras);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed25 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed25 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed25 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_we);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed25 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_we);
		end
		default: begin
			vns_sync_rhs_array_muxed25 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_we);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed26 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed26 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed26 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed26 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			vns_sync_rhs_array_muxed26 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed27 <= 1'd0;
	case (soc_videooverlaysoc_videooverlaysoc_sdram_steerer_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed27 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed27 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed27 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			vns_sync_rhs_array_muxed27 <= ((soc_videooverlaysoc_videooverlaysoc_sdram_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_ready) & soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_is_write);
		end
	endcase
end
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx = vns_xilinxmultiregimpl0_regs1;
assign vns_xilinxasyncresetsynchronizerimpl0 = ((~soc_videooverlaysoc_videooverlaysoc_crg_pll_locked) | soc_videooverlaysoc_videooverlaysoc_crg_rst);
assign vns_xilinxasyncresetsynchronizerimpl1 = ((~soc_videooverlaysoc_videooverlaysoc_crg_pll_locked) | soc_videooverlaysoc_videooverlaysoc_crg_rst);
assign vns_xilinxasyncresetsynchronizerimpl2 = ((~soc_videooverlaysoc_videooverlaysoc_crg_pll_locked) | soc_videooverlaysoc_videooverlaysoc_crg_rst);
assign soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_i = vns_xilinxmultiregimpl1_regs1;
assign soc_videooverlaysoc_hdmi_in0_edid_status = vns_xilinxmultiregimpl2_regs1;
assign soc_videooverlaysoc_hdmi_in0_edid_scl_raw = vns_xilinxmultiregimpl3_regs1;
assign soc_videooverlaysoc_hdmi_in0_edid_sda_raw = vns_xilinxmultiregimpl4_regs1;
assign soc_videooverlaysoc_hdmi_in0_locked = vns_xilinxmultiregimpl5_regs1;
assign vns_xilinxasyncresetsynchronizerimpl3 = (~soc_videooverlaysoc_hdmi_in0_mmcm_locked);
assign vns_xilinxasyncresetsynchronizerimpl4 = (~soc_videooverlaysoc_hdmi_in0_mmcm_locked);
assign vns_xilinxasyncresetsynchronizerimpl5 = (~soc_videooverlaysoc_hdmi_in0_mmcm_locked_o);
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_o = vns_xilinxmultiregimpl6_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_o = vns_xilinxmultiregimpl7_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_o = vns_xilinxmultiregimpl8_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_o = vns_xilinxmultiregimpl9_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_o = vns_xilinxmultiregimpl10_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_status = vns_xilinxmultiregimpl11_regs1;
assign vns_xilinxmultiregimpl11 = {soc_videooverlaysoc_hdmi_in0_s7datacapture0_too_early, soc_videooverlaysoc_hdmi_in0_s7datacapture0_too_late};
assign soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_o = vns_xilinxmultiregimpl12_regs1;
assign soc_videooverlaysoc_hdmi_in0_charsync0_char_synced_status = vns_xilinxmultiregimpl13_regs1;
assign soc_videooverlaysoc_hdmi_in0_charsync0_ctl_pos_status = vns_xilinxmultiregimpl14_regs1;
assign soc_videooverlaysoc_hdmi_in0_wer0_toggle_o = vns_xilinxmultiregimpl15_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_o = vns_xilinxmultiregimpl16_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_o = vns_xilinxmultiregimpl17_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_o = vns_xilinxmultiregimpl18_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_o = vns_xilinxmultiregimpl19_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_o = vns_xilinxmultiregimpl20_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_status = vns_xilinxmultiregimpl21_regs1;
assign vns_xilinxmultiregimpl21 = {soc_videooverlaysoc_hdmi_in0_s7datacapture1_too_early, soc_videooverlaysoc_hdmi_in0_s7datacapture1_too_late};
assign soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_o = vns_xilinxmultiregimpl22_regs1;
assign soc_videooverlaysoc_hdmi_in0_charsync1_char_synced_status = vns_xilinxmultiregimpl23_regs1;
assign soc_videooverlaysoc_hdmi_in0_charsync1_ctl_pos_status = vns_xilinxmultiregimpl24_regs1;
assign soc_videooverlaysoc_hdmi_in0_wer1_toggle_o = vns_xilinxmultiregimpl25_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_o = vns_xilinxmultiregimpl26_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_o = vns_xilinxmultiregimpl27_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_o = vns_xilinxmultiregimpl28_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_o = vns_xilinxmultiregimpl29_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_o = vns_xilinxmultiregimpl30_regs1;
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_status = vns_xilinxmultiregimpl31_regs1;
assign vns_xilinxmultiregimpl31 = {soc_videooverlaysoc_hdmi_in0_s7datacapture2_too_early, soc_videooverlaysoc_hdmi_in0_s7datacapture2_too_late};
assign soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_o = vns_xilinxmultiregimpl32_regs1;
assign soc_videooverlaysoc_hdmi_in0_charsync2_char_synced_status = vns_xilinxmultiregimpl33_regs1;
assign soc_videooverlaysoc_hdmi_in0_charsync2_ctl_pos_status = vns_xilinxmultiregimpl34_regs1;
assign soc_videooverlaysoc_hdmi_in0_wer2_toggle_o = vns_xilinxmultiregimpl35_regs1;
assign soc_videooverlaysoc_hdmi_in0_chansync_status = vns_xilinxmultiregimpl36_regs1;
assign soc_videooverlaysoc_hdmi_in0_decode_terc4_dvimode_bit = vns_xilinxmultiregimpl37_regs1;
assign soc_videooverlaysoc_hdmi_in0_resdetection_hres_status = vns_xilinxmultiregimpl38_regs1;
assign soc_videooverlaysoc_hdmi_in0_resdetection_vres_status = vns_xilinxmultiregimpl39_regs1;
assign soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_i = vns_xilinxmultiregimpl40_regs1;
assign soc_videooverlaysoc_hdmi_in1_edid_scl_raw = vns_xilinxmultiregimpl41_regs1;
assign vns_xilinxmultiregimpl41 = (~hdmi_in1_scl);
assign soc_videooverlaysoc_hdmi_in1_edid_sda_raw = vns_xilinxmultiregimpl42_regs1;
assign soc_videooverlaysoc_hdmi_in1_locked = vns_xilinxmultiregimpl43_regs1;
assign vns_xilinxasyncresetsynchronizerimpl6 = (~soc_videooverlaysoc_hdmi_in1_mmcm_locked);
assign vns_xilinxasyncresetsynchronizerimpl7 = (~soc_videooverlaysoc_hdmi_in1_mmcm_locked);
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_o = vns_xilinxmultiregimpl44_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_o = vns_xilinxmultiregimpl45_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_o = vns_xilinxmultiregimpl46_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_o = vns_xilinxmultiregimpl47_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_o = vns_xilinxmultiregimpl48_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_status = vns_xilinxmultiregimpl49_regs1;
assign vns_xilinxmultiregimpl49 = {soc_videooverlaysoc_hdmi_in1_s7datacapture0_too_early, soc_videooverlaysoc_hdmi_in1_s7datacapture0_too_late};
assign soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_o = vns_xilinxmultiregimpl50_regs1;
assign soc_videooverlaysoc_hdmi_in1_charsync0_char_synced_status = vns_xilinxmultiregimpl51_regs1;
assign soc_videooverlaysoc_hdmi_in1_charsync0_ctl_pos_status = vns_xilinxmultiregimpl52_regs1;
assign soc_videooverlaysoc_hdmi_in1_wer0_toggle_o = vns_xilinxmultiregimpl53_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_o = vns_xilinxmultiregimpl54_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_o = vns_xilinxmultiregimpl55_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_o = vns_xilinxmultiregimpl56_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_o = vns_xilinxmultiregimpl57_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_o = vns_xilinxmultiregimpl58_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_status = vns_xilinxmultiregimpl59_regs1;
assign vns_xilinxmultiregimpl59 = {soc_videooverlaysoc_hdmi_in1_s7datacapture1_too_early, soc_videooverlaysoc_hdmi_in1_s7datacapture1_too_late};
assign soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_o = vns_xilinxmultiregimpl60_regs1;
assign soc_videooverlaysoc_hdmi_in1_charsync1_char_synced_status = vns_xilinxmultiregimpl61_regs1;
assign soc_videooverlaysoc_hdmi_in1_charsync1_ctl_pos_status = vns_xilinxmultiregimpl62_regs1;
assign soc_videooverlaysoc_hdmi_in1_wer1_toggle_o = vns_xilinxmultiregimpl63_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_o = vns_xilinxmultiregimpl64_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_o = vns_xilinxmultiregimpl65_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_o = vns_xilinxmultiregimpl66_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_o = vns_xilinxmultiregimpl67_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_o = vns_xilinxmultiregimpl68_regs1;
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_status = vns_xilinxmultiregimpl69_regs1;
assign vns_xilinxmultiregimpl69 = {soc_videooverlaysoc_hdmi_in1_s7datacapture2_too_early, soc_videooverlaysoc_hdmi_in1_s7datacapture2_too_late};
assign soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_o = vns_xilinxmultiregimpl70_regs1;
assign soc_videooverlaysoc_hdmi_in1_charsync2_char_synced_status = vns_xilinxmultiregimpl71_regs1;
assign soc_videooverlaysoc_hdmi_in1_charsync2_ctl_pos_status = vns_xilinxmultiregimpl72_regs1;
assign soc_videooverlaysoc_hdmi_in1_wer2_toggle_o = vns_xilinxmultiregimpl73_regs1;
assign soc_videooverlaysoc_hdmi_in1_chansync_status = vns_xilinxmultiregimpl74_regs1;
assign soc_videooverlaysoc_hdmi_in1_decode_terc4_dvimode_bit = vns_xilinxmultiregimpl75_regs1;
assign soc_videooverlaysoc_hdmi_in1_resdetection_hres_status = vns_xilinxmultiregimpl76_regs1;
assign soc_videooverlaysoc_hdmi_in1_resdetection_vres_status = vns_xilinxmultiregimpl77_regs1;
assign soc_videooverlaysoc_hdmi_in1_frame_produce_rdomain = vns_xilinxmultiregimpl78_regs1;
assign soc_videooverlaysoc_hdmi_in1_frame_consume_wdomain = vns_xilinxmultiregimpl79_regs1;
assign soc_videooverlaysoc_hdmi_in1_frame_sys_overflow = vns_xilinxmultiregimpl80_regs1;
assign soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_o = vns_xilinxmultiregimpl81_regs1;
assign soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_o = vns_xilinxmultiregimpl82_regs1;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_produce_rdomain = vns_xilinxmultiregimpl83_regs1;
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_consume_wdomain = vns_xilinxmultiregimpl84_regs1;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_produce_rdomain = vns_xilinxmultiregimpl85_regs1;
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_consume_wdomain = vns_xilinxmultiregimpl86_regs1;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_produce_rdomain = vns_xilinxmultiregimpl87_regs1;
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_consume_wdomain = vns_xilinxmultiregimpl88_regs1;
assign soc_videooverlaysoc_hdmi_core_out0_underflow_enable = vns_xilinxmultiregimpl89_regs1;
assign soc_videooverlaysoc_hdmi_core_out0_toggle_o = vns_xilinxmultiregimpl90_regs1;
assign soc_videooverlaysoc_Aksv14 = vns_xilinxmultiregimpl91_regs1;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_valid0 = vns_xilinxmultiregimpl92_regs1;
assign soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_payload_data = vns_xilinxmultiregimpl93_regs1;
assign soc_videooverlaysoc_phy_status = vns_xilinxmultiregimpl94_regs1;
assign soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_o = vns_xilinxmultiregimpl95_regs1;
assign soc_videooverlaysoc_core_mac_ps_crc_error_toggle_o = vns_xilinxmultiregimpl96_regs1;
assign soc_videooverlaysoc_core_mac_tx_cdc_produce_rdomain = vns_xilinxmultiregimpl97_regs1;
assign soc_videooverlaysoc_core_mac_tx_cdc_consume_wdomain = vns_xilinxmultiregimpl98_regs1;
assign soc_videooverlaysoc_core_mac_rx_cdc_produce_rdomain = vns_xilinxmultiregimpl99_regs1;
assign soc_videooverlaysoc_core_mac_rx_cdc_consume_wdomain = vns_xilinxmultiregimpl100_regs1;
assign soc_videooverlaysoc_packet_tx_cdc_produce_rdomain = vns_xilinxmultiregimpl101_regs1;
assign soc_videooverlaysoc_packet_tx_cdc_consume_wdomain = vns_xilinxmultiregimpl102_regs1;
assign soc_videooverlaysoc_packet_rx_cdc_produce_rdomain = vns_xilinxmultiregimpl103_regs1;
assign soc_videooverlaysoc_packet_rx_cdc_consume_wdomain = vns_xilinxmultiregimpl104_regs1;

always @(posedge clk200_clk) begin
	if ((soc_videooverlaysoc_videooverlaysoc_crg_reset_counter != 1'd0)) begin
		soc_videooverlaysoc_videooverlaysoc_crg_reset_counter <= (soc_videooverlaysoc_videooverlaysoc_crg_reset_counter - 1'd1);
	end else begin
		soc_videooverlaysoc_videooverlaysoc_crg_ic_reset <= 1'd0;
	end
	if (clk200_rst) begin
		soc_videooverlaysoc_videooverlaysoc_crg_reset_counter <= 4'd15;
		soc_videooverlaysoc_videooverlaysoc_crg_ic_reset <= 1'd1;
	end
end

always @(posedge eth_clk) begin
	if (soc_videooverlaysoc_phy_counter_ce) begin
		soc_videooverlaysoc_phy_counter <= (soc_videooverlaysoc_phy_counter + 1'd1);
	end
	if (soc_videooverlaysoc_core_mac_ps_preamble_error_o) begin
		soc_videooverlaysoc_core_mac_preamble_errors_status <= (soc_videooverlaysoc_core_mac_preamble_errors_status + 1'd1);
	end
	if (soc_videooverlaysoc_core_mac_ps_crc_error_o) begin
		soc_videooverlaysoc_core_mac_crc_errors_status <= (soc_videooverlaysoc_core_mac_crc_errors_status + 1'd1);
	end
	soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_o_r <= soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_o;
	soc_videooverlaysoc_core_mac_ps_crc_error_toggle_o_r <= soc_videooverlaysoc_core_mac_ps_crc_error_toggle_o;
	soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_binary <= soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_next_binary;
	soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q <= soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_next;
	soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_binary <= soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next_binary;
	soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q <= soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_next;
	case (vns_clockdomainsrenamer1_liteethmac_grant)
		1'd0: begin
			if ((~vns_clockdomainsrenamer1_liteethmac_request[0])) begin
				if (vns_clockdomainsrenamer1_liteethmac_request[1]) begin
					vns_clockdomainsrenamer1_liteethmac_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~vns_clockdomainsrenamer1_liteethmac_request[1])) begin
				if (vns_clockdomainsrenamer1_liteethmac_request[0]) begin
					vns_clockdomainsrenamer1_liteethmac_grant <= 1'd0;
				end
			end
		end
	endcase
	vns_clockdomainsrenamer1_liteethmac_status0_ongoing1 <= ((soc_videooverlaysoc_core_arp_mac_port_sink_valid | vns_clockdomainsrenamer1_liteethmac_status0_ongoing1) & (~vns_clockdomainsrenamer1_liteethmac_status0_last));
	if (vns_clockdomainsrenamer1_liteethmac_status0_last) begin
		vns_clockdomainsrenamer1_liteethmac_status0_first <= 1'd1;
	end else begin
		if ((soc_videooverlaysoc_core_arp_mac_port_sink_valid & soc_videooverlaysoc_core_arp_mac_port_sink_ready)) begin
			vns_clockdomainsrenamer1_liteethmac_status0_first <= 1'd0;
		end
	end
	vns_clockdomainsrenamer1_liteethmac_status1_ongoing1 <= ((soc_videooverlaysoc_core_ip_mac_port_sink_valid | vns_clockdomainsrenamer1_liteethmac_status1_ongoing1) & (~vns_clockdomainsrenamer1_liteethmac_status1_last));
	if (vns_clockdomainsrenamer1_liteethmac_status1_last) begin
		vns_clockdomainsrenamer1_liteethmac_status1_first <= 1'd1;
	end else begin
		if ((soc_videooverlaysoc_core_ip_mac_port_sink_valid & soc_videooverlaysoc_core_ip_mac_port_sink_ready)) begin
			vns_clockdomainsrenamer1_liteethmac_status1_first <= 1'd0;
		end
	end
	if (vns_clockdomainsrenamer1_liteethmac_first) begin
		vns_clockdomainsrenamer1_liteethmac_sel_ongoing <= vns_clockdomainsrenamer1_liteethmac_sel0;
	end
	vns_clockdomainsrenamer1_liteethmac_ongoing1 <= ((soc_videooverlaysoc_core_mac_crossbar_sink_valid | vns_clockdomainsrenamer1_liteethmac_ongoing1) & (~vns_clockdomainsrenamer1_liteethmac_last));
	if (vns_clockdomainsrenamer1_liteethmac_last) begin
		vns_clockdomainsrenamer1_liteethmac_first <= 1'd1;
	end else begin
		if ((soc_videooverlaysoc_core_mac_crossbar_sink_valid & soc_videooverlaysoc_core_mac_crossbar_sink_ready)) begin
			vns_clockdomainsrenamer1_liteethmac_first <= 1'd0;
		end
	end
	if (soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter_reset) begin
		soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter_ce) begin
			soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter <= (soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_mac_liteethmacpacketizer_load) begin
		soc_videooverlaysoc_core_mac_liteethmacpacketizer_header_reg <= soc_videooverlaysoc_core_mac_liteethmacpacketizer_header;
	end else begin
		if (soc_videooverlaysoc_core_mac_liteethmacpacketizer_shift) begin
			soc_videooverlaysoc_core_mac_liteethmacpacketizer_header_reg <= {soc_videooverlaysoc_core_mac_liteethmacpacketizer, soc_videooverlaysoc_core_mac_liteethmacpacketizer_header_reg[111:8]};
		end
	end
	vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_next_state;
	if (soc_videooverlaysoc_core_mac_depacketizer_counter_reset) begin
		soc_videooverlaysoc_core_mac_depacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_mac_depacketizer_counter_ce) begin
			soc_videooverlaysoc_core_mac_depacketizer_counter <= (soc_videooverlaysoc_core_mac_depacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_mac_depacketizer_shift) begin
		soc_videooverlaysoc_core_mac_depacketizer_header_reg <= {soc_videooverlaysoc_core_mac_depacketizer_sink_payload_data, soc_videooverlaysoc_core_mac_depacketizer_header_reg[111:8]};
	end
	if (soc_videooverlaysoc_core_mac_depacketizer_is_el) begin
		soc_videooverlaysoc_core_mac_depacketizer_no_payload <= soc_videooverlaysoc_core_mac_depacketizer_sink_last;
	end
	vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_next_state;
	if (soc_videooverlaysoc_core_arp_tx_counter_reset) begin
		soc_videooverlaysoc_core_arp_tx_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_arp_tx_counter_ce) begin
			soc_videooverlaysoc_core_arp_tx_counter <= (soc_videooverlaysoc_core_arp_tx_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter_reset) begin
		soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter_ce) begin
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter <= (soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_load) begin
		soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header_reg <= soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header;
	end else begin
		if (soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_shift) begin
			soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header_reg <= {soc_videooverlaysoc_core_arp_tx_liteetharppacketizer, soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_header_reg[223:8]};
		end
	end
	vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_state <= vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_next_state;
	vns_clockdomainsrenamer1_liteetharptx_fsm_state <= vns_clockdomainsrenamer1_liteetharptx_fsm_next_state;
	soc_videooverlaysoc_core_arp_valid <= (((((soc_videooverlaysoc_core_arp_depacketizer_source_valid & (soc_videooverlaysoc_core_arp_depacketizer_source_param_hwtype == 1'd1)) & (soc_videooverlaysoc_core_arp_depacketizer_source_param_proto == 12'd2048)) & (soc_videooverlaysoc_core_arp_depacketizer_source_param_hwsize == 3'd6)) & (soc_videooverlaysoc_core_arp_depacketizer_source_param_protosize == 3'd4)) & (soc_videooverlaysoc_core_arp_depacketizer_source_param_target_ip == 28'd167774978));
	if (soc_videooverlaysoc_core_arp_depacketizer_counter_reset) begin
		soc_videooverlaysoc_core_arp_depacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_arp_depacketizer_counter_ce) begin
			soc_videooverlaysoc_core_arp_depacketizer_counter <= (soc_videooverlaysoc_core_arp_depacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_arp_depacketizer_shift) begin
		soc_videooverlaysoc_core_arp_depacketizer_header_reg <= {soc_videooverlaysoc_core_arp_depacketizer_sink_payload_data, soc_videooverlaysoc_core_arp_depacketizer_header_reg[223:8]};
	end
	if (soc_videooverlaysoc_core_arp_depacketizer_is_el) begin
		soc_videooverlaysoc_core_arp_depacketizer_no_payload <= soc_videooverlaysoc_core_arp_depacketizer_sink_last;
	end
	vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_state <= vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_next_state;
	vns_clockdomainsrenamer1_liteetharprx_fsm_state <= vns_clockdomainsrenamer1_liteetharprx_fsm_next_state;
	if (soc_videooverlaysoc_core_arp_table_request_pending_clr) begin
		soc_videooverlaysoc_core_arp_table_request_pending <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_arp_table_request_pending_set) begin
			soc_videooverlaysoc_core_arp_table_request_pending <= 1'd1;
		end
	end
	if (soc_videooverlaysoc_core_arp_table_request_ip_address_reset) begin
		soc_videooverlaysoc_core_arp_table_request_ip_address <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_arp_table_request_ip_address_update) begin
			soc_videooverlaysoc_core_arp_table_request_ip_address <= soc_videooverlaysoc_core_arp_table_request_payload_ip_address;
		end
	end
	if (soc_videooverlaysoc_core_arp_table_request_counter_reset) begin
		soc_videooverlaysoc_core_arp_table_request_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_arp_table_request_counter_ce) begin
			soc_videooverlaysoc_core_arp_table_request_counter <= (soc_videooverlaysoc_core_arp_table_request_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_arp_table_update) begin
		soc_videooverlaysoc_core_arp_table_cached_valid <= 1'd1;
		soc_videooverlaysoc_core_arp_table_cached_ip_address <= soc_videooverlaysoc_core_arp_table_sink_payload_ip_address;
		soc_videooverlaysoc_core_arp_table_cached_mac_address <= soc_videooverlaysoc_core_arp_table_sink_payload_mac_address;
	end else begin
		if (soc_videooverlaysoc_core_arp_table_cached_timer_done) begin
			soc_videooverlaysoc_core_arp_table_cached_valid <= 1'd0;
		end
	end
	if (soc_videooverlaysoc_core_arp_table_request_timer_wait) begin
		if ((~soc_videooverlaysoc_core_arp_table_request_timer_done)) begin
			soc_videooverlaysoc_core_arp_table_request_timer_count <= (soc_videooverlaysoc_core_arp_table_request_timer_count - 1'd1);
		end
	end else begin
		soc_videooverlaysoc_core_arp_table_request_timer_count <= 23'd5000000;
	end
	if (soc_videooverlaysoc_core_arp_table_cached_timer_wait) begin
		if ((~soc_videooverlaysoc_core_arp_table_cached_timer_done)) begin
			soc_videooverlaysoc_core_arp_table_cached_timer_count <= (soc_videooverlaysoc_core_arp_table_cached_timer_count - 1'd1);
		end
	end else begin
		soc_videooverlaysoc_core_arp_table_cached_timer_count <= 29'd500000000;
	end
	vns_clockdomainsrenamer1_state1 <= vns_clockdomainsrenamer1_next_state1;
	if (soc_videooverlaysoc_core_arp_table_response_valid) begin
		soc_videooverlaysoc_core_ip_tx_target_mac <= soc_videooverlaysoc_core_arp_table_response_payload_mac_address;
	end
	if (soc_videooverlaysoc_core_ip_tx_ce) begin
		if ((~soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next0 <= {soc_videooverlaysoc_core_ip_tx_liteethipv4checksum0, (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next0[15:0] + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next0[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next1 <= {soc_videooverlaysoc_core_ip_tx_liteethipv4checksum1, (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next1[15:0] + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next1[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next2 <= {soc_videooverlaysoc_core_ip_tx_liteethipv4checksum2, (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next2[15:0] + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next2[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next3 <= {soc_videooverlaysoc_core_ip_tx_liteethipv4checksum3, (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next3[15:0] + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next3[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next4 <= {soc_videooverlaysoc_core_ip_tx_liteethipv4checksum4, (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next4[15:0] + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next4[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next5 <= {soc_videooverlaysoc_core_ip_tx_liteethipv4checksum5, (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next5[15:0] + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next5[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next6 <= {soc_videooverlaysoc_core_ip_tx_liteethipv4checksum6, (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next6[15:0] + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next6[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next7 <= {soc_videooverlaysoc_core_ip_tx_liteethipv4checksum7, (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next7[15:0] + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next7[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_r_next8 <= {soc_videooverlaysoc_core_ip_tx_liteethipv4checksum8, (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next8[15:0] + soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_s_next8[16])};
		end
		if (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_counter_ce) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_counter <= (soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_ip_tx_reset) begin
		soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_counter <= 4'd0;
	end
	if (soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter_reset) begin
		soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter_ce) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter <= (soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_load) begin
		soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header_reg <= soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header;
	end else begin
		if (soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_shift) begin
			soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header_reg <= {soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer, soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_header_reg[159:8]};
		end
	end
	vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_state <= vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_next_state;
	vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_state <= vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_next_state;
	soc_videooverlaysoc_core_ip_rx_valid <= ((((soc_videooverlaysoc_core_ip_rx_depacketizer_source_valid & (soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_target_ip == 28'd167774978)) & (soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_version == 3'd4)) & (soc_videooverlaysoc_core_ip_rx_depacketizer_source_param_ihl == 3'd5)) & (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_value == 1'd0));
	if (soc_videooverlaysoc_core_ip_rx_depacketizer_counter_reset) begin
		soc_videooverlaysoc_core_ip_rx_depacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_ip_rx_depacketizer_counter_ce) begin
			soc_videooverlaysoc_core_ip_rx_depacketizer_counter <= (soc_videooverlaysoc_core_ip_rx_depacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_ip_rx_depacketizer_shift) begin
		soc_videooverlaysoc_core_ip_rx_depacketizer_header_reg <= {soc_videooverlaysoc_core_ip_rx_depacketizer_sink_payload_data, soc_videooverlaysoc_core_ip_rx_depacketizer_header_reg[159:8]};
	end
	if (soc_videooverlaysoc_core_ip_rx_depacketizer_is_el) begin
		soc_videooverlaysoc_core_ip_rx_depacketizer_no_payload <= soc_videooverlaysoc_core_ip_rx_depacketizer_sink_last;
	end
	vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_state <= vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_next_state;
	if (soc_videooverlaysoc_core_ip_rx_ce) begin
		if ((~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next0 <= {soc_videooverlaysoc_core_ip_rx_liteethipv4checksum0, (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next0[15:0] + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next0[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next1 <= {soc_videooverlaysoc_core_ip_rx_liteethipv4checksum1, (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next1[15:0] + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next1[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next2 <= {soc_videooverlaysoc_core_ip_rx_liteethipv4checksum2, (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next2[15:0] + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next2[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next3 <= {soc_videooverlaysoc_core_ip_rx_liteethipv4checksum3, (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next3[15:0] + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next3[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next4 <= {soc_videooverlaysoc_core_ip_rx_liteethipv4checksum4, (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next4[15:0] + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next4[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next5 <= {soc_videooverlaysoc_core_ip_rx_liteethipv4checksum5, (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next5[15:0] + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next5[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next6 <= {soc_videooverlaysoc_core_ip_rx_liteethipv4checksum6, (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next6[15:0] + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next6[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next7 <= {soc_videooverlaysoc_core_ip_rx_liteethipv4checksum7, (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next7[15:0] + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next7[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next8 <= {soc_videooverlaysoc_core_ip_rx_liteethipv4checksum8, (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next8[15:0] + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next8[16])};
		end
		if ((~soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_done)) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_r_next9 <= {soc_videooverlaysoc_core_ip_rx_liteethipv4checksum9, (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next9[15:0] + soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_s_next9[16])};
		end
		if (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_counter_ce) begin
			soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_counter <= (soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_ip_rx_reset) begin
		soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_counter <= 4'd0;
	end
	vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_state <= vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_next_state;
	case (vns_clockdomainsrenamer1_liteethip_grant)
		1'd0: begin
			if ((~vns_clockdomainsrenamer1_liteethip_request[0])) begin
				if (vns_clockdomainsrenamer1_liteethip_request[1]) begin
					vns_clockdomainsrenamer1_liteethip_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~vns_clockdomainsrenamer1_liteethip_request[1])) begin
				if (vns_clockdomainsrenamer1_liteethip_request[0]) begin
					vns_clockdomainsrenamer1_liteethip_grant <= 1'd0;
				end
			end
		end
	endcase
	vns_clockdomainsrenamer1_liteethip_status0_ongoing1 <= ((soc_videooverlaysoc_core_icmp_ip_port_sink_valid | vns_clockdomainsrenamer1_liteethip_status0_ongoing1) & (~vns_clockdomainsrenamer1_liteethip_status0_last));
	if (vns_clockdomainsrenamer1_liteethip_status0_last) begin
		vns_clockdomainsrenamer1_liteethip_status0_first <= 1'd1;
	end else begin
		if ((soc_videooverlaysoc_core_icmp_ip_port_sink_valid & soc_videooverlaysoc_core_icmp_ip_port_sink_ready)) begin
			vns_clockdomainsrenamer1_liteethip_status0_first <= 1'd0;
		end
	end
	vns_clockdomainsrenamer1_liteethip_status1_ongoing1 <= ((soc_videooverlaysoc_core_ip_port_sink_valid | vns_clockdomainsrenamer1_liteethip_status1_ongoing1) & (~vns_clockdomainsrenamer1_liteethip_status1_last));
	if (vns_clockdomainsrenamer1_liteethip_status1_last) begin
		vns_clockdomainsrenamer1_liteethip_status1_first <= 1'd1;
	end else begin
		if ((soc_videooverlaysoc_core_ip_port_sink_valid & soc_videooverlaysoc_core_ip_port_sink_ready)) begin
			vns_clockdomainsrenamer1_liteethip_status1_first <= 1'd0;
		end
	end
	if (vns_clockdomainsrenamer1_liteethip_first) begin
		vns_clockdomainsrenamer1_liteethip_sel_ongoing <= vns_clockdomainsrenamer1_liteethip_sel0;
	end
	vns_clockdomainsrenamer1_liteethip_ongoing1 <= ((soc_videooverlaysoc_core_ip_crossbar_sink_valid | vns_clockdomainsrenamer1_liteethip_ongoing1) & (~vns_clockdomainsrenamer1_liteethip_last));
	if (vns_clockdomainsrenamer1_liteethip_last) begin
		vns_clockdomainsrenamer1_liteethip_first <= 1'd1;
	end else begin
		if ((soc_videooverlaysoc_core_ip_crossbar_sink_valid & soc_videooverlaysoc_core_ip_crossbar_sink_ready)) begin
			vns_clockdomainsrenamer1_liteethip_first <= 1'd0;
		end
	end
	if (soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter_reset) begin
		soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter_ce) begin
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter <= (soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_load) begin
		soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header_reg <= soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header;
	end else begin
		if (soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_shift) begin
			soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header_reg <= {soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer, soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_header_reg[63:8]};
		end
	end
	vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_state <= vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_next_state;
	vns_clockdomainsrenamer1_liteethicmptx_fsm_state <= vns_clockdomainsrenamer1_liteethicmptx_fsm_next_state;
	soc_videooverlaysoc_core_icmp_rx_valid <= (soc_videooverlaysoc_core_icmp_rx_depacketizer_source_valid & (soc_videooverlaysoc_core_icmp_rx_sink_sink_param_protocol == 1'd1));
	if (soc_videooverlaysoc_core_icmp_rx_depacketizer_counter_reset) begin
		soc_videooverlaysoc_core_icmp_rx_depacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_icmp_rx_depacketizer_counter_ce) begin
			soc_videooverlaysoc_core_icmp_rx_depacketizer_counter <= (soc_videooverlaysoc_core_icmp_rx_depacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_icmp_rx_depacketizer_shift) begin
		soc_videooverlaysoc_core_icmp_rx_depacketizer_header_reg <= {soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_payload_data, soc_videooverlaysoc_core_icmp_rx_depacketizer_header_reg[63:8]};
	end
	if (soc_videooverlaysoc_core_icmp_rx_depacketizer_is_el) begin
		soc_videooverlaysoc_core_icmp_rx_depacketizer_no_payload <= soc_videooverlaysoc_core_icmp_rx_depacketizer_sink_last;
	end
	vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_state <= vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_next_state;
	vns_clockdomainsrenamer1_liteethicmprx_fsm_state <= vns_clockdomainsrenamer1_liteethicmprx_fsm_next_state;
	if (soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_re) begin
		soc_videooverlaysoc_core_icmp_echo_buffer_readable <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_core_icmp_echo_buffer_re) begin
			soc_videooverlaysoc_core_icmp_echo_buffer_readable <= 1'd0;
		end
	end
	if (((soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_we & soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_writable) & (~soc_videooverlaysoc_core_icmp_echo_buffer_replace))) begin
		soc_videooverlaysoc_core_icmp_echo_buffer_produce <= (soc_videooverlaysoc_core_icmp_echo_buffer_produce + 1'd1);
	end
	if (soc_videooverlaysoc_core_icmp_echo_buffer_do_read) begin
		soc_videooverlaysoc_core_icmp_echo_buffer_consume <= (soc_videooverlaysoc_core_icmp_echo_buffer_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_we & soc_videooverlaysoc_core_icmp_echo_buffer_syncfifo_writable) & (~soc_videooverlaysoc_core_icmp_echo_buffer_replace))) begin
		if ((~soc_videooverlaysoc_core_icmp_echo_buffer_do_read)) begin
			soc_videooverlaysoc_core_icmp_echo_buffer_level0 <= (soc_videooverlaysoc_core_icmp_echo_buffer_level0 + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_core_icmp_echo_buffer_do_read) begin
			soc_videooverlaysoc_core_icmp_echo_buffer_level0 <= (soc_videooverlaysoc_core_icmp_echo_buffer_level0 - 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_tx_liteethudppacketizer_counter_reset) begin
		soc_videooverlaysoc_core_tx_liteethudppacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_tx_liteethudppacketizer_counter_ce) begin
			soc_videooverlaysoc_core_tx_liteethudppacketizer_counter <= (soc_videooverlaysoc_core_tx_liteethudppacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_tx_liteethudppacketizer_load) begin
		soc_videooverlaysoc_core_tx_liteethudppacketizer_header_reg <= soc_videooverlaysoc_core_tx_liteethudppacketizer_header;
	end else begin
		if (soc_videooverlaysoc_core_tx_liteethudppacketizer_shift) begin
			soc_videooverlaysoc_core_tx_liteethudppacketizer_header_reg <= {soc_videooverlaysoc_core_tx_liteethudppacketizer, soc_videooverlaysoc_core_tx_liteethudppacketizer_header_reg[63:8]};
		end
	end
	vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_state <= vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_next_state;
	vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_state <= vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_next_state;
	soc_videooverlaysoc_core_valid <= (soc_videooverlaysoc_core_depacketizer_source_valid & (soc_videooverlaysoc_core_sink_sink_param_protocol == 5'd17));
	if (soc_videooverlaysoc_core_depacketizer_counter_reset) begin
		soc_videooverlaysoc_core_depacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_depacketizer_counter_ce) begin
			soc_videooverlaysoc_core_depacketizer_counter <= (soc_videooverlaysoc_core_depacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_depacketizer_shift) begin
		soc_videooverlaysoc_core_depacketizer_header_reg <= {soc_videooverlaysoc_core_depacketizer_sink_payload_data, soc_videooverlaysoc_core_depacketizer_header_reg[63:8]};
	end
	if (soc_videooverlaysoc_core_depacketizer_is_el) begin
		soc_videooverlaysoc_core_depacketizer_no_payload <= soc_videooverlaysoc_core_depacketizer_sink_last;
	end
	vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_state <= vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_next_state;
	vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_state <= vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_next_state;
	soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_binary <= soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next_binary;
	soc_videooverlaysoc_packet_tx_cdc_graycounter1_q <= soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_next;
	if ((soc_videooverlaysoc_packet_tx_converter_converter_source_valid & soc_videooverlaysoc_packet_tx_converter_converter_source_ready)) begin
		if (soc_videooverlaysoc_packet_tx_converter_converter_last) begin
			soc_videooverlaysoc_packet_tx_converter_converter_mux <= 1'd0;
		end else begin
			soc_videooverlaysoc_packet_tx_converter_converter_mux <= (soc_videooverlaysoc_packet_tx_converter_converter_mux + 1'd1);
		end
	end
	soc_videooverlaysoc_packet_rx_converter_source_param_src_port <= soc_videooverlaysoc_packet_rx_converter_sink_param_src_port;
	soc_videooverlaysoc_packet_rx_converter_source_param_dst_port <= soc_videooverlaysoc_packet_rx_converter_sink_param_dst_port;
	soc_videooverlaysoc_packet_rx_converter_source_param_ip_address <= soc_videooverlaysoc_packet_rx_converter_sink_param_ip_address;
	soc_videooverlaysoc_packet_rx_converter_source_param_length <= soc_videooverlaysoc_packet_rx_converter_sink_param_length;
	if (soc_videooverlaysoc_packet_rx_converter_converter_source_ready) begin
		soc_videooverlaysoc_packet_rx_converter_converter_strobe_all <= 1'd0;
	end
	if (soc_videooverlaysoc_packet_rx_converter_converter_load_part) begin
		if (((soc_videooverlaysoc_packet_rx_converter_converter_demux == 2'd3) | soc_videooverlaysoc_packet_rx_converter_converter_sink_last)) begin
			soc_videooverlaysoc_packet_rx_converter_converter_demux <= 1'd0;
			soc_videooverlaysoc_packet_rx_converter_converter_strobe_all <= 1'd1;
		end else begin
			soc_videooverlaysoc_packet_rx_converter_converter_demux <= (soc_videooverlaysoc_packet_rx_converter_converter_demux + 1'd1);
		end
	end
	if ((soc_videooverlaysoc_packet_rx_converter_converter_source_valid & soc_videooverlaysoc_packet_rx_converter_converter_source_ready)) begin
		if ((soc_videooverlaysoc_packet_rx_converter_converter_sink_valid & soc_videooverlaysoc_packet_rx_converter_converter_sink_ready)) begin
			soc_videooverlaysoc_packet_rx_converter_converter_source_first <= soc_videooverlaysoc_packet_rx_converter_converter_sink_first;
			soc_videooverlaysoc_packet_rx_converter_converter_source_last <= soc_videooverlaysoc_packet_rx_converter_converter_sink_last;
		end else begin
			soc_videooverlaysoc_packet_rx_converter_converter_source_first <= 1'd0;
			soc_videooverlaysoc_packet_rx_converter_converter_source_last <= 1'd0;
		end
	end else begin
		if ((soc_videooverlaysoc_packet_rx_converter_converter_sink_valid & soc_videooverlaysoc_packet_rx_converter_converter_sink_ready)) begin
			soc_videooverlaysoc_packet_rx_converter_converter_source_first <= (soc_videooverlaysoc_packet_rx_converter_converter_sink_first | soc_videooverlaysoc_packet_rx_converter_converter_source_first);
			soc_videooverlaysoc_packet_rx_converter_converter_source_last <= (soc_videooverlaysoc_packet_rx_converter_converter_sink_last | soc_videooverlaysoc_packet_rx_converter_converter_source_last);
		end
	end
	if (soc_videooverlaysoc_packet_rx_converter_converter_load_part) begin
		case (soc_videooverlaysoc_packet_rx_converter_converter_demux)
			1'd0: begin
				soc_videooverlaysoc_packet_rx_converter_converter_source_payload_data[8:0] <= soc_videooverlaysoc_packet_rx_converter_converter_sink_payload_data;
			end
			1'd1: begin
				soc_videooverlaysoc_packet_rx_converter_converter_source_payload_data[17:9] <= soc_videooverlaysoc_packet_rx_converter_converter_sink_payload_data;
			end
			2'd2: begin
				soc_videooverlaysoc_packet_rx_converter_converter_source_payload_data[26:18] <= soc_videooverlaysoc_packet_rx_converter_converter_sink_payload_data;
			end
			2'd3: begin
				soc_videooverlaysoc_packet_rx_converter_converter_source_payload_data[35:27] <= soc_videooverlaysoc_packet_rx_converter_converter_sink_payload_data;
			end
		endcase
	end
	if (soc_videooverlaysoc_packet_rx_converter_converter_load_part) begin
		soc_videooverlaysoc_packet_rx_converter_converter_source_payload_valid_token_count <= (soc_videooverlaysoc_packet_rx_converter_converter_demux + 1'd1);
	end
	soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_binary <= soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_next_binary;
	soc_videooverlaysoc_packet_rx_cdc_graycounter0_q <= soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_next;
	if (eth_rst) begin
		soc_videooverlaysoc_phy_counter <= 9'd0;
		soc_videooverlaysoc_core_mac_preamble_errors_status <= 32'd0;
		soc_videooverlaysoc_core_mac_crc_errors_status <= 32'd0;
		soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q <= 7'd0;
		soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q_binary <= 7'd0;
		soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q <= 7'd0;
		soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q_binary <= 7'd0;
		soc_videooverlaysoc_core_mac_liteethmacpacketizer_counter <= 4'd0;
		soc_videooverlaysoc_core_mac_depacketizer_counter <= 4'd0;
		soc_videooverlaysoc_core_mac_depacketizer_no_payload <= 1'd0;
		soc_videooverlaysoc_core_arp_tx_liteetharppacketizer_counter <= 5'd0;
		soc_videooverlaysoc_core_arp_depacketizer_counter <= 5'd0;
		soc_videooverlaysoc_core_arp_depacketizer_no_payload <= 1'd0;
		soc_videooverlaysoc_core_arp_table_request_pending <= 1'd0;
		soc_videooverlaysoc_core_arp_table_request_timer_count <= 23'd5000000;
		soc_videooverlaysoc_core_arp_table_request_counter <= 3'd0;
		soc_videooverlaysoc_core_arp_table_cached_valid <= 1'd0;
		soc_videooverlaysoc_core_arp_table_cached_timer_count <= 29'd500000000;
		soc_videooverlaysoc_core_ip_tx_liteethipv4checksum_counter <= 4'd0;
		soc_videooverlaysoc_core_ip_tx_liteethipv4packetizer_counter <= 5'd0;
		soc_videooverlaysoc_core_ip_rx_depacketizer_counter <= 5'd0;
		soc_videooverlaysoc_core_ip_rx_depacketizer_no_payload <= 1'd0;
		soc_videooverlaysoc_core_ip_rx_liteethipv4checksum_counter <= 4'd0;
		soc_videooverlaysoc_core_icmp_tx_liteethicmppacketizer_counter <= 3'd0;
		soc_videooverlaysoc_core_icmp_rx_depacketizer_counter <= 3'd0;
		soc_videooverlaysoc_core_icmp_rx_depacketizer_no_payload <= 1'd0;
		soc_videooverlaysoc_core_icmp_echo_buffer_readable <= 1'd0;
		soc_videooverlaysoc_core_icmp_echo_buffer_level0 <= 8'd0;
		soc_videooverlaysoc_core_icmp_echo_buffer_produce <= 7'd0;
		soc_videooverlaysoc_core_icmp_echo_buffer_consume <= 7'd0;
		soc_videooverlaysoc_core_tx_liteethudppacketizer_counter <= 3'd0;
		soc_videooverlaysoc_core_depacketizer_counter <= 3'd0;
		soc_videooverlaysoc_core_depacketizer_no_payload <= 1'd0;
		soc_videooverlaysoc_packet_tx_cdc_graycounter1_q <= 3'd0;
		soc_videooverlaysoc_packet_tx_cdc_graycounter1_q_binary <= 3'd0;
		soc_videooverlaysoc_packet_tx_converter_converter_mux <= 2'd0;
		soc_videooverlaysoc_packet_rx_converter_source_param_src_port <= 16'd0;
		soc_videooverlaysoc_packet_rx_converter_source_param_dst_port <= 16'd0;
		soc_videooverlaysoc_packet_rx_converter_source_param_ip_address <= 32'd0;
		soc_videooverlaysoc_packet_rx_converter_source_param_length <= 16'd0;
		soc_videooverlaysoc_packet_rx_converter_converter_source_first <= 1'd0;
		soc_videooverlaysoc_packet_rx_converter_converter_source_last <= 1'd0;
		soc_videooverlaysoc_packet_rx_converter_converter_source_payload_data <= 36'd0;
		soc_videooverlaysoc_packet_rx_converter_converter_source_payload_valid_token_count <= 3'd0;
		soc_videooverlaysoc_packet_rx_converter_converter_demux <= 2'd0;
		soc_videooverlaysoc_packet_rx_converter_converter_strobe_all <= 1'd0;
		soc_videooverlaysoc_packet_rx_cdc_graycounter0_q <= 3'd0;
		soc_videooverlaysoc_packet_rx_cdc_graycounter0_q_binary <= 3'd0;
		vns_clockdomainsrenamer1_liteethmac_grant <= 1'd0;
		vns_clockdomainsrenamer1_liteethmac_status0_first <= 1'd1;
		vns_clockdomainsrenamer1_liteethmac_status0_ongoing1 <= 1'd0;
		vns_clockdomainsrenamer1_liteethmac_status1_first <= 1'd1;
		vns_clockdomainsrenamer1_liteethmac_status1_ongoing1 <= 1'd0;
		vns_clockdomainsrenamer1_liteethmac_first <= 1'd1;
		vns_clockdomainsrenamer1_liteethmac_ongoing1 <= 1'd0;
		vns_clockdomainsrenamer1_liteethmac_sel_ongoing <= 2'd0;
		vns_clockdomainsrenamer1_liteethmac_liteethmacpacketizer_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethmac_liteethmacdepacketizer_state <= 2'd0;
		vns_clockdomainsrenamer1_liteetharptx_liteetharppacketizer_state <= 2'd0;
		vns_clockdomainsrenamer1_liteetharptx_fsm_state <= 1'd0;
		vns_clockdomainsrenamer1_liteetharprx_liteetharpdepacketizer_state <= 2'd0;
		vns_clockdomainsrenamer1_liteetharprx_fsm_state <= 2'd0;
		vns_clockdomainsrenamer1_state1 <= 3'd0;
		vns_clockdomainsrenamer1_liteethip_liteethiptx_liteethipv4packetizer_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethip_liteethiptx_fsm_state <= 3'd0;
		vns_clockdomainsrenamer1_liteethip_liteethiprx_liteethipv4depacketizer_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethip_liteethiprx_fsm_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethip_grant <= 1'd0;
		vns_clockdomainsrenamer1_liteethip_status0_first <= 1'd1;
		vns_clockdomainsrenamer1_liteethip_status0_ongoing1 <= 1'd0;
		vns_clockdomainsrenamer1_liteethip_status1_first <= 1'd1;
		vns_clockdomainsrenamer1_liteethip_status1_ongoing1 <= 1'd0;
		vns_clockdomainsrenamer1_liteethip_first <= 1'd1;
		vns_clockdomainsrenamer1_liteethip_ongoing1 <= 1'd0;
		vns_clockdomainsrenamer1_liteethip_sel_ongoing <= 2'd0;
		vns_clockdomainsrenamer1_liteethicmptx_liteethicmppacketizer_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethicmptx_fsm_state <= 1'd0;
		vns_clockdomainsrenamer1_liteethicmprx_liteethicmpdepacketizer_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethicmprx_fsm_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethudp_liteethudptx_liteethudppacketizer_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethudp_liteethudptx_fsm_state <= 1'd0;
		vns_clockdomainsrenamer1_liteethudp_liteethudprx_liteethudpdepacketizer_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethudp_liteethudprx_fsm_state <= 2'd0;
	end
	vns_xilinxmultiregimpl94_regs0 <= soc_videooverlaysoc_phy_data_r;
	vns_xilinxmultiregimpl94_regs1 <= vns_xilinxmultiregimpl94_regs0;
	vns_xilinxmultiregimpl95_regs0 <= soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_i;
	vns_xilinxmultiregimpl95_regs1 <= vns_xilinxmultiregimpl95_regs0;
	vns_xilinxmultiregimpl96_regs0 <= soc_videooverlaysoc_core_mac_ps_crc_error_toggle_i;
	vns_xilinxmultiregimpl96_regs1 <= vns_xilinxmultiregimpl96_regs0;
	vns_xilinxmultiregimpl98_regs0 <= soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q;
	vns_xilinxmultiregimpl98_regs1 <= vns_xilinxmultiregimpl98_regs0;
	vns_xilinxmultiregimpl99_regs0 <= soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q;
	vns_xilinxmultiregimpl99_regs1 <= vns_xilinxmultiregimpl99_regs0;
	vns_xilinxmultiregimpl101_regs0 <= soc_videooverlaysoc_packet_tx_cdc_graycounter0_q;
	vns_xilinxmultiregimpl101_regs1 <= vns_xilinxmultiregimpl101_regs0;
	vns_xilinxmultiregimpl104_regs0 <= soc_videooverlaysoc_packet_rx_cdc_graycounter1_q;
	vns_xilinxmultiregimpl104_regs1 <= vns_xilinxmultiregimpl104_regs0;
end

always @(posedge eth_rx_clk) begin
	soc_videooverlaysoc_phy_liteethphyrmiirx_crs_dv <= rmii_eth_crs_dv;
	soc_videooverlaysoc_phy_liteethphyrmiirx_crs_dv_d <= soc_videooverlaysoc_phy_liteethphyrmiirx_crs_dv;
	soc_videooverlaysoc_phy_liteethphyrmiirx_rx_data <= rmii_eth_rx_data;
	if (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_ready) begin
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_strobe_all <= 1'd0;
	end
	if (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_load_part) begin
		if (((soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_demux == 2'd3) | soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_last)) begin
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_demux <= 1'd0;
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_strobe_all <= 1'd1;
		end else begin
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_demux <= (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_demux + 1'd1);
		end
	end
	if ((soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_valid & soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_ready)) begin
		if ((soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_valid & soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_ready)) begin
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_first <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_first;
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_last <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_last;
		end else begin
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_first <= 1'd0;
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_last <= 1'd0;
		end
	end else begin
		if ((soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_valid & soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_ready)) begin
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_first <= (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_first | soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_first);
			soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_last <= (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_last | soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_last);
		end
	end
	if (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_load_part) begin
		case (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_demux)
			1'd0: begin
				soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_data[1:0] <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_payload_data;
			end
			1'd1: begin
				soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_data[3:2] <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_payload_data;
			end
			2'd2: begin
				soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_data[5:4] <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_payload_data;
			end
			2'd3: begin
				soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_data[7:6] <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_sink_payload_data;
			end
		endcase
	end
	if (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_load_part) begin
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_valid_token_count <= (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_demux + 1'd1);
	end
	if (soc_videooverlaysoc_phy_liteethphyrmiirx_converter_reset) begin
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_first <= 1'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_last <= 1'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_data <= 8'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_valid_token_count <= 3'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_demux <= 2'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_strobe_all <= 1'd0;
	end
	vns_clockdomainsrenamer0_state1 <= vns_clockdomainsrenamer0_next_state1;
	vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_next_state;
	if (soc_videooverlaysoc_core_mac_crc32_checker_crc_ce) begin
		soc_videooverlaysoc_core_mac_crc32_checker_crc_reg <= soc_videooverlaysoc_core_mac_crc32_checker_crc_next;
	end
	if (soc_videooverlaysoc_core_mac_crc32_checker_crc_reset) begin
		soc_videooverlaysoc_core_mac_crc32_checker_crc_reg <= 32'd4294967295;
	end
	if (((soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_we & soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_writable) & (~soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_replace))) begin
		if ((soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_produce == 3'd4)) begin
			soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_produce <= 1'd0;
		end else begin
			soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_produce <= (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_produce + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_do_read) begin
		if ((soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_consume == 3'd4)) begin
			soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_consume <= 1'd0;
		end else begin
			soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_consume <= (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_consume + 1'd1);
		end
	end
	if (((soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_we & soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_syncfifo_writable) & (~soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_replace))) begin
		if ((~soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_do_read)) begin
			soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_level <= (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_do_read) begin
			soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_level <= (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_mac_crc32_checker_fifo_reset) begin
		soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_level <= 3'd0;
		soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_produce <= 3'd0;
		soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_consume <= 3'd0;
	end
	vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_state <= vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_next_state;
	if (soc_videooverlaysoc_core_mac_ps_preamble_error_i) begin
		soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_i <= (~soc_videooverlaysoc_core_mac_ps_preamble_error_toggle_i);
	end
	if (soc_videooverlaysoc_core_mac_ps_crc_error_i) begin
		soc_videooverlaysoc_core_mac_ps_crc_error_toggle_i <= (~soc_videooverlaysoc_core_mac_ps_crc_error_toggle_i);
	end
	soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_binary <= soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_next_binary;
	soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q <= soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_next;
	if (eth_rx_rst) begin
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_first <= 1'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_last <= 1'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_data <= 8'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_source_payload_valid_token_count <= 3'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_demux <= 2'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_converter_converter_strobe_all <= 1'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_crs_dv <= 1'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_crs_dv_d <= 1'd0;
		soc_videooverlaysoc_phy_liteethphyrmiirx_rx_data <= 2'd0;
		soc_videooverlaysoc_core_mac_crc32_checker_crc_reg <= 32'd4294967295;
		soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_level <= 3'd0;
		soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_produce <= 3'd0;
		soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_consume <= 3'd0;
		soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q <= 7'd0;
		soc_videooverlaysoc_core_mac_rx_cdc_graycounter0_q_binary <= 7'd0;
		vns_clockdomainsrenamer0_state1 <= 1'd0;
		vns_clockdomainsrenamer1_liteethmac_liteethmacpreamblechecker_state <= 1'd0;
		vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32checker_state <= 2'd0;
	end
	vns_xilinxmultiregimpl92_regs0 <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_valid1;
	vns_xilinxmultiregimpl92_regs1 <= vns_xilinxmultiregimpl92_regs0;
	vns_xilinxmultiregimpl93_regs0 <= soc_videooverlaysoc_phy_liteethphyrmiirx_converter_sink_data;
	vns_xilinxmultiregimpl93_regs1 <= vns_xilinxmultiregimpl93_regs0;
	vns_xilinxmultiregimpl100_regs0 <= soc_videooverlaysoc_core_mac_rx_cdc_graycounter1_q;
	vns_xilinxmultiregimpl100_regs1 <= vns_xilinxmultiregimpl100_regs0;
end

always @(posedge eth_tx_clk) begin
	rmii_eth_tx_en <= soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_valid;
	rmii_eth_tx_data <= soc_videooverlaysoc_phy_liteethphyrmiitx_converter_source_payload_data;
	if ((soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_valid & soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_source_ready)) begin
		if (soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_last) begin
			soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_mux <= 1'd0;
		end else begin
			soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_mux <= (soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_mux + 1'd1);
		end
	end
	if (soc_videooverlaysoc_core_mac_tx_gap_inserter_counter_reset) begin
		soc_videooverlaysoc_core_mac_tx_gap_inserter_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_mac_tx_gap_inserter_counter_ce) begin
			soc_videooverlaysoc_core_mac_tx_gap_inserter_counter <= (soc_videooverlaysoc_core_mac_tx_gap_inserter_counter + 1'd1);
		end
	end
	vns_clockdomainsrenamer1_liteethmac_liteethmacgap_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacgap_next_state;
	if (soc_videooverlaysoc_core_mac_preamble_inserter_clr_cnt) begin
		soc_videooverlaysoc_core_mac_preamble_inserter_cnt <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_mac_preamble_inserter_inc_cnt) begin
			soc_videooverlaysoc_core_mac_preamble_inserter_cnt <= (soc_videooverlaysoc_core_mac_preamble_inserter_cnt + 1'd1);
		end
	end
	vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_next_state;
	if (soc_videooverlaysoc_core_mac_crc32_inserter_is_ongoing0) begin
		soc_videooverlaysoc_core_mac_crc32_inserter_cnt <= 2'd3;
	end else begin
		if ((soc_videooverlaysoc_core_mac_crc32_inserter_is_ongoing1 & (~soc_videooverlaysoc_core_mac_crc32_inserter_cnt_done))) begin
			soc_videooverlaysoc_core_mac_crc32_inserter_cnt <= (soc_videooverlaysoc_core_mac_crc32_inserter_cnt - soc_videooverlaysoc_core_mac_crc32_inserter_source_ready);
		end
	end
	if (soc_videooverlaysoc_core_mac_crc32_inserter_ce) begin
		soc_videooverlaysoc_core_mac_crc32_inserter_reg <= soc_videooverlaysoc_core_mac_crc32_inserter_next;
	end
	if (soc_videooverlaysoc_core_mac_crc32_inserter_reset) begin
		soc_videooverlaysoc_core_mac_crc32_inserter_reg <= 32'd4294967295;
	end
	vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_state <= vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_next_state;
	if (soc_videooverlaysoc_core_mac_padding_inserter_counter_reset) begin
		soc_videooverlaysoc_core_mac_padding_inserter_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_core_mac_padding_inserter_counter_ce) begin
			soc_videooverlaysoc_core_mac_padding_inserter_counter <= (soc_videooverlaysoc_core_mac_padding_inserter_counter + 1'd1);
		end
	end
	vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_state <= vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_next_state;
	soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_binary <= soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next_binary;
	soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q <= soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_next;
	if (eth_tx_rst) begin
		soc_videooverlaysoc_phy_liteethphyrmiitx_converter_converter_mux <= 2'd0;
		soc_videooverlaysoc_core_mac_crc32_inserter_reg <= 32'd4294967295;
		soc_videooverlaysoc_core_mac_crc32_inserter_cnt <= 2'd3;
		soc_videooverlaysoc_core_mac_padding_inserter_counter <= 16'd1;
		soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q <= 7'd0;
		soc_videooverlaysoc_core_mac_tx_cdc_graycounter1_q_binary <= 7'd0;
		vns_clockdomainsrenamer1_liteethmac_liteethmacgap_state <= 1'd0;
		vns_clockdomainsrenamer1_liteethmac_liteethmacpreambleinserter_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethmac_liteethmaccrc32inserter_state <= 2'd0;
		vns_clockdomainsrenamer1_liteethmac_liteethmacpaddinginserter_state <= 1'd0;
	end
	vns_xilinxmultiregimpl97_regs0 <= soc_videooverlaysoc_core_mac_tx_cdc_graycounter0_q;
	vns_xilinxmultiregimpl97_regs1 <= vns_xilinxmultiregimpl97_regs0;
end

always @(posedge etherbone_clk) begin
	soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_binary <= soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_next_binary;
	soc_videooverlaysoc_packet_tx_cdc_graycounter0_q <= soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_next;
	soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_binary <= soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next_binary;
	soc_videooverlaysoc_packet_rx_cdc_graycounter1_q <= soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_next;
	if (etherbone_rst) begin
		soc_videooverlaysoc_packet_tx_cdc_graycounter0_q <= 3'd0;
		soc_videooverlaysoc_packet_tx_cdc_graycounter0_q_binary <= 3'd0;
		soc_videooverlaysoc_packet_rx_cdc_graycounter1_q <= 3'd0;
		soc_videooverlaysoc_packet_rx_cdc_graycounter1_q_binary <= 3'd0;
	end
	vns_xilinxmultiregimpl102_regs0 <= soc_videooverlaysoc_packet_tx_cdc_graycounter1_q;
	vns_xilinxmultiregimpl102_regs1 <= vns_xilinxmultiregimpl102_regs0;
	vns_xilinxmultiregimpl103_regs0 <= soc_videooverlaysoc_packet_rx_cdc_graycounter0_q;
	vns_xilinxmultiregimpl103_regs1 <= vns_xilinxmultiregimpl103_regs0;
end

always @(posedge hdmi_in0_data0_cap_read_clk) begin
	soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst_read <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst;
	soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_rd <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr;
	if ((soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rdpointer == 3'd7)) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rdpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rdpointer <= (soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rdpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rdpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_rd[9:0];
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_rd[19:10];
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_rd[29:20];
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_rd[39:30];
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_rd[49:40];
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_rd[59:50];
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_rd[69:60];
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_rd[79:70];
		end
	endcase
	if (hdmi_in0_data0_cap_read_rst) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst_read <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge hdmi_in0_data0_cap_write_clk) begin
	soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst_write <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst;
	if ((soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_wrpointer == 4'd9)) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_wrpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_wrpointer <= (soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_wrpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_wrpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr[7:0] <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr[15:8] <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr[23:16] <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr[31:24] <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr[39:32] <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr[47:40] <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr[55:48] <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr[63:56] <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
		end
		4'd8: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr[71:64] <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
		end
		4'd9: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_storage_wr[79:72] <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_i;
		end
	endcase
	if (hdmi_in0_data0_cap_write_rst) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_rst_write <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge hdmi_in0_data1_cap_read_clk) begin
	soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst_read <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst;
	soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_rd <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr;
	if ((soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rdpointer == 3'd7)) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rdpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rdpointer <= (soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rdpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rdpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_rd[9:0];
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_rd[19:10];
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_rd[29:20];
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_rd[39:30];
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_rd[49:40];
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_rd[59:50];
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_rd[69:60];
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_rd[79:70];
		end
	endcase
	if (hdmi_in0_data1_cap_read_rst) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst_read <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge hdmi_in0_data1_cap_write_clk) begin
	soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst_write <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst;
	if ((soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_wrpointer == 4'd9)) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_wrpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_wrpointer <= (soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_wrpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_wrpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr[7:0] <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr[15:8] <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr[23:16] <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr[31:24] <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr[39:32] <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr[47:40] <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr[55:48] <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr[63:56] <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
		end
		4'd8: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr[71:64] <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
		end
		4'd9: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_storage_wr[79:72] <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_i;
		end
	endcase
	if (hdmi_in0_data1_cap_write_rst) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_rst_write <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge hdmi_in0_data2_cap_read_clk) begin
	soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst_read <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst;
	soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_rd <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr;
	if ((soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rdpointer == 3'd7)) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rdpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rdpointer <= (soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rdpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rdpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_rd[9:0];
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_rd[19:10];
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_rd[29:20];
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_rd[39:30];
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_rd[49:40];
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_rd[59:50];
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_rd[69:60];
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_rd[79:70];
		end
	endcase
	if (hdmi_in0_data2_cap_read_rst) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst_read <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge hdmi_in0_data2_cap_write_clk) begin
	soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst_write <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst;
	if ((soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_wrpointer == 4'd9)) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_wrpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_wrpointer <= (soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_wrpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_wrpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr[7:0] <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr[15:8] <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr[23:16] <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr[31:24] <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr[39:32] <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr[47:40] <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr[55:48] <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr[63:56] <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
		end
		4'd8: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr[71:64] <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
		end
		4'd9: begin
			soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_storage_wr[79:72] <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_i;
		end
	endcase
	if (hdmi_in0_data2_cap_write_rst) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_rst_write <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge hdmi_in0_freq_fmeter_clk) begin
	soc_videooverlaysoc_hdmi_in0_freq_q_binary <= soc_videooverlaysoc_hdmi_in0_freq_q_next_binary;
	soc_videooverlaysoc_hdmi_in0_freq_q <= soc_videooverlaysoc_hdmi_in0_freq_q_next;
end

always @(posedge hdmi_in0_pix_clk) begin
	soc_videooverlaysoc_hdmi_in0_charsync0_raw_data1 <= soc_videooverlaysoc_hdmi_in0_charsync0_raw_data;
	soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd0;
	if (((((soc_videooverlaysoc_hdmi_in0_charsync0_raw[9:0] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[9:0] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[9:0] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[9:0] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 1'd0;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync0_raw[10:1] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[10:1] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[10:1] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[10:1] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 1'd1;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync0_raw[11:2] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[11:2] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[11:2] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[11:2] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 2'd2;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync0_raw[12:3] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[12:3] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[12:3] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[12:3] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 2'd3;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync0_raw[13:4] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[13:4] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[13:4] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[13:4] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 3'd4;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync0_raw[14:5] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[14:5] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[14:5] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[14:5] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 3'd5;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync0_raw[15:6] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[15:6] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[15:6] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[15:6] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 3'd6;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync0_raw[16:7] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[16:7] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[16:7] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[16:7] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 3'd7;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync0_raw[17:8] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[17:8] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[17:8] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[17:8] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 4'd8;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync0_raw[18:9] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[18:9] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[18:9] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync0_raw[18:9] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in0_charsync0_found_control & (soc_videooverlaysoc_hdmi_in0_charsync0_control_position == soc_videooverlaysoc_hdmi_in0_charsync0_previous_control_position))) begin
		if ((soc_videooverlaysoc_hdmi_in0_charsync0_control_counter == 3'd7)) begin
			soc_videooverlaysoc_hdmi_in0_charsync0_control_counter <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_charsync0_synced <= 1'd1;
			soc_videooverlaysoc_hdmi_in0_charsync0_word_sel <= soc_videooverlaysoc_hdmi_in0_charsync0_control_position;
		end else begin
			soc_videooverlaysoc_hdmi_in0_charsync0_control_counter <= (soc_videooverlaysoc_hdmi_in0_charsync0_control_counter + 1'd1);
		end
	end else begin
		soc_videooverlaysoc_hdmi_in0_charsync0_control_counter <= 1'd0;
	end
	soc_videooverlaysoc_hdmi_in0_charsync0_previous_control_position <= soc_videooverlaysoc_hdmi_in0_charsync0_control_position;
	soc_videooverlaysoc_hdmi_in0_charsync0_data <= (soc_videooverlaysoc_hdmi_in0_charsync0_raw >>> soc_videooverlaysoc_hdmi_in0_charsync0_word_sel);
	soc_videooverlaysoc_hdmi_in0_wer0_data_r <= soc_videooverlaysoc_hdmi_in0_wer0_data[8:0];
	soc_videooverlaysoc_hdmi_in0_wer0_transition_count <= (((((((soc_videooverlaysoc_hdmi_in0_wer0_transitions[0] + soc_videooverlaysoc_hdmi_in0_wer0_transitions[1]) + soc_videooverlaysoc_hdmi_in0_wer0_transitions[2]) + soc_videooverlaysoc_hdmi_in0_wer0_transitions[3]) + soc_videooverlaysoc_hdmi_in0_wer0_transitions[4]) + soc_videooverlaysoc_hdmi_in0_wer0_transitions[5]) + soc_videooverlaysoc_hdmi_in0_wer0_transitions[6]) + soc_videooverlaysoc_hdmi_in0_wer0_transitions[7]);
	soc_videooverlaysoc_hdmi_in0_wer0_is_control <= ((((soc_videooverlaysoc_hdmi_in0_wer0_data_r == 10'd852) | (soc_videooverlaysoc_hdmi_in0_wer0_data_r == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_wer0_data_r == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_wer0_data_r == 10'd683));
	soc_videooverlaysoc_hdmi_in0_wer0_is_error <= ((soc_videooverlaysoc_hdmi_in0_wer0_transition_count > 3'd4) & (~soc_videooverlaysoc_hdmi_in0_wer0_is_control));
	{soc_videooverlaysoc_hdmi_in0_wer0_period_done, soc_videooverlaysoc_hdmi_in0_wer0_period_counter} <= (soc_videooverlaysoc_hdmi_in0_wer0_period_counter + 1'd1);
	soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_r_updated <= soc_videooverlaysoc_hdmi_in0_wer0_period_done;
	if (soc_videooverlaysoc_hdmi_in0_wer0_period_done) begin
		soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_r <= soc_videooverlaysoc_hdmi_in0_wer0_wer_counter;
		soc_videooverlaysoc_hdmi_in0_wer0_wer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in0_wer0_is_error) begin
			soc_videooverlaysoc_hdmi_in0_wer0_wer_counter <= (soc_videooverlaysoc_hdmi_in0_wer0_wer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in0_wer0_i) begin
		soc_videooverlaysoc_hdmi_in0_wer0_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_wer0_toggle_i);
	end
	soc_videooverlaysoc_hdmi_in0_decoding0_output_de <= 1'd1;
	if ((soc_videooverlaysoc_hdmi_in0_decoding0_input == 10'd852)) begin
		soc_videooverlaysoc_hdmi_in0_decoding0_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding0_output_c <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decoding0_input == 8'd171)) begin
		soc_videooverlaysoc_hdmi_in0_decoding0_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding0_output_c <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decoding0_input == 9'd340)) begin
		soc_videooverlaysoc_hdmi_in0_decoding0_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding0_output_c <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decoding0_input == 10'd683)) begin
		soc_videooverlaysoc_hdmi_in0_decoding0_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding0_output_c <= 2'd3;
	end
	soc_videooverlaysoc_hdmi_in0_decoding0_output_raw <= soc_videooverlaysoc_hdmi_in0_decoding0_input;
	soc_videooverlaysoc_hdmi_in0_decoding0_output_d[0] <= (soc_videooverlaysoc_hdmi_in0_decoding0_input[0] ^ soc_videooverlaysoc_hdmi_in0_decoding0_input[9]);
	soc_videooverlaysoc_hdmi_in0_decoding0_output_d[1] <= ((soc_videooverlaysoc_hdmi_in0_decoding0_input[1] ^ soc_videooverlaysoc_hdmi_in0_decoding0_input[0]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding0_output_d[2] <= ((soc_videooverlaysoc_hdmi_in0_decoding0_input[2] ^ soc_videooverlaysoc_hdmi_in0_decoding0_input[1]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding0_output_d[3] <= ((soc_videooverlaysoc_hdmi_in0_decoding0_input[3] ^ soc_videooverlaysoc_hdmi_in0_decoding0_input[2]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding0_output_d[4] <= ((soc_videooverlaysoc_hdmi_in0_decoding0_input[4] ^ soc_videooverlaysoc_hdmi_in0_decoding0_input[3]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding0_output_d[5] <= ((soc_videooverlaysoc_hdmi_in0_decoding0_input[5] ^ soc_videooverlaysoc_hdmi_in0_decoding0_input[4]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding0_output_d[6] <= ((soc_videooverlaysoc_hdmi_in0_decoding0_input[6] ^ soc_videooverlaysoc_hdmi_in0_decoding0_input[5]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding0_output_d[7] <= ((soc_videooverlaysoc_hdmi_in0_decoding0_input[7] ^ soc_videooverlaysoc_hdmi_in0_decoding0_input[6]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding0_valid_o <= soc_videooverlaysoc_hdmi_in0_decoding0_valid_i;
	soc_videooverlaysoc_hdmi_in0_charsync1_raw_data1 <= soc_videooverlaysoc_hdmi_in0_charsync1_raw_data;
	soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd0;
	if (((((soc_videooverlaysoc_hdmi_in0_charsync1_raw[9:0] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[9:0] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[9:0] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[9:0] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 1'd0;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync1_raw[10:1] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[10:1] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[10:1] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[10:1] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 1'd1;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync1_raw[11:2] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[11:2] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[11:2] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[11:2] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 2'd2;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync1_raw[12:3] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[12:3] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[12:3] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[12:3] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 2'd3;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync1_raw[13:4] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[13:4] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[13:4] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[13:4] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 3'd4;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync1_raw[14:5] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[14:5] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[14:5] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[14:5] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 3'd5;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync1_raw[15:6] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[15:6] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[15:6] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[15:6] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 3'd6;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync1_raw[16:7] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[16:7] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[16:7] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[16:7] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 3'd7;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync1_raw[17:8] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[17:8] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[17:8] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[17:8] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 4'd8;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync1_raw[18:9] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[18:9] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[18:9] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync1_raw[18:9] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in0_charsync1_found_control & (soc_videooverlaysoc_hdmi_in0_charsync1_control_position == soc_videooverlaysoc_hdmi_in0_charsync1_previous_control_position))) begin
		if ((soc_videooverlaysoc_hdmi_in0_charsync1_control_counter == 3'd7)) begin
			soc_videooverlaysoc_hdmi_in0_charsync1_control_counter <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_charsync1_synced <= 1'd1;
			soc_videooverlaysoc_hdmi_in0_charsync1_word_sel <= soc_videooverlaysoc_hdmi_in0_charsync1_control_position;
		end else begin
			soc_videooverlaysoc_hdmi_in0_charsync1_control_counter <= (soc_videooverlaysoc_hdmi_in0_charsync1_control_counter + 1'd1);
		end
	end else begin
		soc_videooverlaysoc_hdmi_in0_charsync1_control_counter <= 1'd0;
	end
	soc_videooverlaysoc_hdmi_in0_charsync1_previous_control_position <= soc_videooverlaysoc_hdmi_in0_charsync1_control_position;
	soc_videooverlaysoc_hdmi_in0_charsync1_data <= (soc_videooverlaysoc_hdmi_in0_charsync1_raw >>> soc_videooverlaysoc_hdmi_in0_charsync1_word_sel);
	soc_videooverlaysoc_hdmi_in0_wer1_data_r <= soc_videooverlaysoc_hdmi_in0_wer1_data[8:0];
	soc_videooverlaysoc_hdmi_in0_wer1_transition_count <= (((((((soc_videooverlaysoc_hdmi_in0_wer1_transitions[0] + soc_videooverlaysoc_hdmi_in0_wer1_transitions[1]) + soc_videooverlaysoc_hdmi_in0_wer1_transitions[2]) + soc_videooverlaysoc_hdmi_in0_wer1_transitions[3]) + soc_videooverlaysoc_hdmi_in0_wer1_transitions[4]) + soc_videooverlaysoc_hdmi_in0_wer1_transitions[5]) + soc_videooverlaysoc_hdmi_in0_wer1_transitions[6]) + soc_videooverlaysoc_hdmi_in0_wer1_transitions[7]);
	soc_videooverlaysoc_hdmi_in0_wer1_is_control <= ((((soc_videooverlaysoc_hdmi_in0_wer1_data_r == 10'd852) | (soc_videooverlaysoc_hdmi_in0_wer1_data_r == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_wer1_data_r == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_wer1_data_r == 10'd683));
	soc_videooverlaysoc_hdmi_in0_wer1_is_error <= ((soc_videooverlaysoc_hdmi_in0_wer1_transition_count > 3'd4) & (~soc_videooverlaysoc_hdmi_in0_wer1_is_control));
	{soc_videooverlaysoc_hdmi_in0_wer1_period_done, soc_videooverlaysoc_hdmi_in0_wer1_period_counter} <= (soc_videooverlaysoc_hdmi_in0_wer1_period_counter + 1'd1);
	soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_r_updated <= soc_videooverlaysoc_hdmi_in0_wer1_period_done;
	if (soc_videooverlaysoc_hdmi_in0_wer1_period_done) begin
		soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_r <= soc_videooverlaysoc_hdmi_in0_wer1_wer_counter;
		soc_videooverlaysoc_hdmi_in0_wer1_wer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in0_wer1_is_error) begin
			soc_videooverlaysoc_hdmi_in0_wer1_wer_counter <= (soc_videooverlaysoc_hdmi_in0_wer1_wer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in0_wer1_i) begin
		soc_videooverlaysoc_hdmi_in0_wer1_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_wer1_toggle_i);
	end
	soc_videooverlaysoc_hdmi_in0_decoding1_output_de <= 1'd1;
	if ((soc_videooverlaysoc_hdmi_in0_decoding1_input == 10'd852)) begin
		soc_videooverlaysoc_hdmi_in0_decoding1_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding1_output_c <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decoding1_input == 8'd171)) begin
		soc_videooverlaysoc_hdmi_in0_decoding1_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding1_output_c <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decoding1_input == 9'd340)) begin
		soc_videooverlaysoc_hdmi_in0_decoding1_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding1_output_c <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decoding1_input == 10'd683)) begin
		soc_videooverlaysoc_hdmi_in0_decoding1_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding1_output_c <= 2'd3;
	end
	soc_videooverlaysoc_hdmi_in0_decoding1_output_raw <= soc_videooverlaysoc_hdmi_in0_decoding1_input;
	soc_videooverlaysoc_hdmi_in0_decoding1_output_d[0] <= (soc_videooverlaysoc_hdmi_in0_decoding1_input[0] ^ soc_videooverlaysoc_hdmi_in0_decoding1_input[9]);
	soc_videooverlaysoc_hdmi_in0_decoding1_output_d[1] <= ((soc_videooverlaysoc_hdmi_in0_decoding1_input[1] ^ soc_videooverlaysoc_hdmi_in0_decoding1_input[0]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding1_output_d[2] <= ((soc_videooverlaysoc_hdmi_in0_decoding1_input[2] ^ soc_videooverlaysoc_hdmi_in0_decoding1_input[1]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding1_output_d[3] <= ((soc_videooverlaysoc_hdmi_in0_decoding1_input[3] ^ soc_videooverlaysoc_hdmi_in0_decoding1_input[2]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding1_output_d[4] <= ((soc_videooverlaysoc_hdmi_in0_decoding1_input[4] ^ soc_videooverlaysoc_hdmi_in0_decoding1_input[3]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding1_output_d[5] <= ((soc_videooverlaysoc_hdmi_in0_decoding1_input[5] ^ soc_videooverlaysoc_hdmi_in0_decoding1_input[4]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding1_output_d[6] <= ((soc_videooverlaysoc_hdmi_in0_decoding1_input[6] ^ soc_videooverlaysoc_hdmi_in0_decoding1_input[5]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding1_output_d[7] <= ((soc_videooverlaysoc_hdmi_in0_decoding1_input[7] ^ soc_videooverlaysoc_hdmi_in0_decoding1_input[6]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding1_valid_o <= soc_videooverlaysoc_hdmi_in0_decoding1_valid_i;
	soc_videooverlaysoc_hdmi_in0_charsync2_raw_data1 <= soc_videooverlaysoc_hdmi_in0_charsync2_raw_data;
	soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd0;
	if (((((soc_videooverlaysoc_hdmi_in0_charsync2_raw[9:0] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[9:0] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[9:0] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[9:0] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 1'd0;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync2_raw[10:1] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[10:1] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[10:1] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[10:1] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 1'd1;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync2_raw[11:2] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[11:2] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[11:2] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[11:2] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 2'd2;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync2_raw[12:3] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[12:3] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[12:3] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[12:3] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 2'd3;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync2_raw[13:4] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[13:4] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[13:4] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[13:4] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 3'd4;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync2_raw[14:5] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[14:5] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[14:5] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[14:5] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 3'd5;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync2_raw[15:6] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[15:6] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[15:6] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[15:6] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 3'd6;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync2_raw[16:7] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[16:7] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[16:7] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[16:7] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 3'd7;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync2_raw[17:8] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[17:8] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[17:8] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[17:8] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 4'd8;
	end
	if (((((soc_videooverlaysoc_hdmi_in0_charsync2_raw[18:9] == 10'd852) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[18:9] == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[18:9] == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_charsync2_raw[18:9] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in0_charsync2_found_control & (soc_videooverlaysoc_hdmi_in0_charsync2_control_position == soc_videooverlaysoc_hdmi_in0_charsync2_previous_control_position))) begin
		if ((soc_videooverlaysoc_hdmi_in0_charsync2_control_counter == 3'd7)) begin
			soc_videooverlaysoc_hdmi_in0_charsync2_control_counter <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_charsync2_synced <= 1'd1;
			soc_videooverlaysoc_hdmi_in0_charsync2_word_sel <= soc_videooverlaysoc_hdmi_in0_charsync2_control_position;
		end else begin
			soc_videooverlaysoc_hdmi_in0_charsync2_control_counter <= (soc_videooverlaysoc_hdmi_in0_charsync2_control_counter + 1'd1);
		end
	end else begin
		soc_videooverlaysoc_hdmi_in0_charsync2_control_counter <= 1'd0;
	end
	soc_videooverlaysoc_hdmi_in0_charsync2_previous_control_position <= soc_videooverlaysoc_hdmi_in0_charsync2_control_position;
	soc_videooverlaysoc_hdmi_in0_charsync2_data <= (soc_videooverlaysoc_hdmi_in0_charsync2_raw >>> soc_videooverlaysoc_hdmi_in0_charsync2_word_sel);
	soc_videooverlaysoc_hdmi_in0_wer2_data_r <= soc_videooverlaysoc_hdmi_in0_wer2_data[8:0];
	soc_videooverlaysoc_hdmi_in0_wer2_transition_count <= (((((((soc_videooverlaysoc_hdmi_in0_wer2_transitions[0] + soc_videooverlaysoc_hdmi_in0_wer2_transitions[1]) + soc_videooverlaysoc_hdmi_in0_wer2_transitions[2]) + soc_videooverlaysoc_hdmi_in0_wer2_transitions[3]) + soc_videooverlaysoc_hdmi_in0_wer2_transitions[4]) + soc_videooverlaysoc_hdmi_in0_wer2_transitions[5]) + soc_videooverlaysoc_hdmi_in0_wer2_transitions[6]) + soc_videooverlaysoc_hdmi_in0_wer2_transitions[7]);
	soc_videooverlaysoc_hdmi_in0_wer2_is_control <= ((((soc_videooverlaysoc_hdmi_in0_wer2_data_r == 10'd852) | (soc_videooverlaysoc_hdmi_in0_wer2_data_r == 8'd171)) | (soc_videooverlaysoc_hdmi_in0_wer2_data_r == 9'd340)) | (soc_videooverlaysoc_hdmi_in0_wer2_data_r == 10'd683));
	soc_videooverlaysoc_hdmi_in0_wer2_is_error <= ((soc_videooverlaysoc_hdmi_in0_wer2_transition_count > 3'd4) & (~soc_videooverlaysoc_hdmi_in0_wer2_is_control));
	{soc_videooverlaysoc_hdmi_in0_wer2_period_done, soc_videooverlaysoc_hdmi_in0_wer2_period_counter} <= (soc_videooverlaysoc_hdmi_in0_wer2_period_counter + 1'd1);
	soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_r_updated <= soc_videooverlaysoc_hdmi_in0_wer2_period_done;
	if (soc_videooverlaysoc_hdmi_in0_wer2_period_done) begin
		soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_r <= soc_videooverlaysoc_hdmi_in0_wer2_wer_counter;
		soc_videooverlaysoc_hdmi_in0_wer2_wer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in0_wer2_is_error) begin
			soc_videooverlaysoc_hdmi_in0_wer2_wer_counter <= (soc_videooverlaysoc_hdmi_in0_wer2_wer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in0_wer2_i) begin
		soc_videooverlaysoc_hdmi_in0_wer2_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_wer2_toggle_i);
	end
	soc_videooverlaysoc_hdmi_in0_decoding2_output_de <= 1'd1;
	if ((soc_videooverlaysoc_hdmi_in0_decoding2_input == 10'd852)) begin
		soc_videooverlaysoc_hdmi_in0_decoding2_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding2_output_c <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decoding2_input == 8'd171)) begin
		soc_videooverlaysoc_hdmi_in0_decoding2_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding2_output_c <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decoding2_input == 9'd340)) begin
		soc_videooverlaysoc_hdmi_in0_decoding2_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding2_output_c <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decoding2_input == 10'd683)) begin
		soc_videooverlaysoc_hdmi_in0_decoding2_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding2_output_c <= 2'd3;
	end
	soc_videooverlaysoc_hdmi_in0_decoding2_output_raw <= soc_videooverlaysoc_hdmi_in0_decoding2_input;
	soc_videooverlaysoc_hdmi_in0_decoding2_output_d[0] <= (soc_videooverlaysoc_hdmi_in0_decoding2_input[0] ^ soc_videooverlaysoc_hdmi_in0_decoding2_input[9]);
	soc_videooverlaysoc_hdmi_in0_decoding2_output_d[1] <= ((soc_videooverlaysoc_hdmi_in0_decoding2_input[1] ^ soc_videooverlaysoc_hdmi_in0_decoding2_input[0]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding2_output_d[2] <= ((soc_videooverlaysoc_hdmi_in0_decoding2_input[2] ^ soc_videooverlaysoc_hdmi_in0_decoding2_input[1]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding2_output_d[3] <= ((soc_videooverlaysoc_hdmi_in0_decoding2_input[3] ^ soc_videooverlaysoc_hdmi_in0_decoding2_input[2]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding2_output_d[4] <= ((soc_videooverlaysoc_hdmi_in0_decoding2_input[4] ^ soc_videooverlaysoc_hdmi_in0_decoding2_input[3]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding2_output_d[5] <= ((soc_videooverlaysoc_hdmi_in0_decoding2_input[5] ^ soc_videooverlaysoc_hdmi_in0_decoding2_input[4]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding2_output_d[6] <= ((soc_videooverlaysoc_hdmi_in0_decoding2_input[6] ^ soc_videooverlaysoc_hdmi_in0_decoding2_input[5]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding2_output_d[7] <= ((soc_videooverlaysoc_hdmi_in0_decoding2_input[7] ^ soc_videooverlaysoc_hdmi_in0_decoding2_input[6]) ^ (~soc_videooverlaysoc_hdmi_in0_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in0_decoding2_valid_o <= soc_videooverlaysoc_hdmi_in0_decoding2_valid_i;
	if ((~soc_videooverlaysoc_hdmi_in0_chansync_valid_i)) begin
		soc_videooverlaysoc_hdmi_in0_chansync_chan_synced <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in0_chansync_some_control) begin
			if (soc_videooverlaysoc_hdmi_in0_chansync_all_control) begin
				soc_videooverlaysoc_hdmi_in0_chansync_chan_synced <= 1'd1;
			end else begin
				soc_videooverlaysoc_hdmi_in0_chansync_chan_synced <= 1'd0;
			end
		end
	end
	soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_produce <= (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_produce + 1'd1);
	if (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_re) begin
		soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_consume <= (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_consume + 1'd1);
	end
	soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_produce <= (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_produce + 1'd1);
	if (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_re) begin
		soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_consume <= (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_consume + 1'd1);
	end
	soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_produce <= (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_produce + 1'd1);
	if (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_re) begin
		soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_consume <= (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_consume + 1'd1);
	end
	soc_videooverlaysoc_hdmi_in0_decode_terc4_de_r <= soc_videooverlaysoc_hdmi_in0_decode_terc4_data_in0_de;
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd668)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd611)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd740)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd738)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 2'd3;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 9'd369)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 3'd4;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 9'd286)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 3'd5;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 9'd398)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 3'd6;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 9'd316)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 3'd7;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd716)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd8;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 9'd313)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 9'd412)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd10;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd710)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd11;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd654)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd12;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd625)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd13;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 9'd355)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd14;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd707)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd15;
	end
	if (soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_valid_in) begin
		if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd852)) begin
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd1;
		end else begin
			if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 8'd171)) begin
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c <= 1'd1;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd1;
			end else begin
				if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 9'd340)) begin
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c <= 2'd2;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd1;
				end else begin
					if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd683)) begin
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c <= 2'd3;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd1;
					end else begin
						if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 9'd307)) begin
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c <= 1'd0;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd1;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd0;
						end else begin
							if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_data_in_raw == 10'd716)) begin
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd1;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd0;
							end else begin
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd1;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd0;
							end
						end
					end
				end
			end
		end
	end else begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd668)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd611)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd740)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd738)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 2'd3;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 9'd369)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 3'd4;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 9'd286)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 3'd5;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 9'd398)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 3'd6;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 9'd316)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 3'd7;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd716)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd8;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 9'd313)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 9'd412)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd10;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd710)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd11;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd654)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd12;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd625)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd13;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 9'd355)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd14;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd707)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd15;
	end
	if (soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_valid_in) begin
		if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd852)) begin
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd1;
		end else begin
			if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 8'd171)) begin
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c <= 1'd1;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd1;
			end else begin
				if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 9'd340)) begin
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c <= 2'd2;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd1;
				end else begin
					if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 10'd683)) begin
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c <= 2'd3;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd1;
					end else begin
						if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 9'd307)) begin
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c <= 1'd0;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd1;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd1;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd0;
						end else begin
							if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_data_in_raw == 9'd307)) begin
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd1;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd1;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd0;
							end else begin
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd1;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd0;
							end
						end
					end
				end
			end
		end
	end else begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd668)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd611)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd740)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd738)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 2'd3;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 9'd369)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 3'd4;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 9'd286)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 3'd5;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 9'd398)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 3'd6;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 9'd316)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 3'd7;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd716)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd8;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 9'd313)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 9'd412)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd10;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd710)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd11;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd654)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd12;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd625)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd13;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 9'd355)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd14;
	end
	if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd707)) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd15;
	end
	if (soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_valid_in) begin
		if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd852)) begin
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd1;
		end else begin
			if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 8'd171)) begin
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c <= 1'd1;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd1;
			end else begin
				if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 9'd340)) begin
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c <= 2'd2;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd1;
				end else begin
					if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd683)) begin
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c <= 2'd3;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd1;
					end else begin
						if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 9'd307)) begin
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c <= 1'd0;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd1;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
							soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd0;
						end else begin
							if ((soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_data_in_raw == 10'd716)) begin
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd1;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd0;
							end else begin
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd1;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd0;
							end
						end
					end
				end
			end
		end
	end else begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd0;
	end
	vns_clockdomainsrenamer0_state0 <= vns_clockdomainsrenamer0_next_state0;
	soc_videooverlaysoc_hdmi_in0_syncpol_valid_o <= soc_videooverlaysoc_hdmi_in0_syncpol_valid_i;
	soc_videooverlaysoc_hdmi_in0_syncpol_r <= soc_videooverlaysoc_hdmi_in0_syncpol_data_in2_d;
	soc_videooverlaysoc_hdmi_in0_syncpol_g <= soc_videooverlaysoc_hdmi_in0_syncpol_data_in1_d;
	soc_videooverlaysoc_hdmi_in0_syncpol_b <= soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_d;
	soc_videooverlaysoc_hdmi_in0_syncpol_de_r <= soc_videooverlaysoc_hdmi_in0_syncpol_de_int;
	if (soc_videooverlaysoc_hdmi_in0_syncpol_de_rising) begin
		soc_videooverlaysoc_hdmi_in0_syncpol_c_polarity <= soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_c;
		soc_videooverlaysoc_hdmi_in0_syncpol_c_out <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in0_syncpol_c_out <= (soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_c ^ soc_videooverlaysoc_hdmi_in0_syncpol_c_polarity);
	end
	soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s0 <= soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_raw;
	soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s1 <= soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_d;
	soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s2 <= soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_c;
	soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s3 <= soc_videooverlaysoc_hdmi_in0_data0_timingdelay_sink_de;
	soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s0 <= soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_raw;
	soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s1 <= soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_d;
	soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s2 <= soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_c;
	soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s3 <= soc_videooverlaysoc_hdmi_in0_data1_timingdelay_sink_de;
	soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s0 <= soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_raw;
	soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s1 <= soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_d;
	soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s2 <= soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_c;
	soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s3 <= soc_videooverlaysoc_hdmi_in0_data2_timingdelay_sink_de;
	soc_videooverlaysoc_hdmi_in0_resdetection_de_r <= soc_videooverlaysoc_hdmi_in0_resdetection_de;
	if ((soc_videooverlaysoc_hdmi_in0_resdetection_valid_i & soc_videooverlaysoc_hdmi_in0_resdetection_de)) begin
		soc_videooverlaysoc_hdmi_in0_resdetection_hcounter <= (soc_videooverlaysoc_hdmi_in0_resdetection_hcounter + 1'd1);
	end else begin
		soc_videooverlaysoc_hdmi_in0_resdetection_hcounter <= 1'd0;
	end
	if (soc_videooverlaysoc_hdmi_in0_resdetection_valid_i) begin
		if (soc_videooverlaysoc_hdmi_in0_resdetection_pn_de) begin
			soc_videooverlaysoc_hdmi_in0_resdetection_hcounter_st <= soc_videooverlaysoc_hdmi_in0_resdetection_hcounter;
		end
	end else begin
		soc_videooverlaysoc_hdmi_in0_resdetection_hcounter_st <= 1'd0;
	end
	soc_videooverlaysoc_hdmi_in0_resdetection_vsync_r <= soc_videooverlaysoc_hdmi_in0_resdetection_vsync;
	if ((soc_videooverlaysoc_hdmi_in0_resdetection_valid_i & soc_videooverlaysoc_hdmi_in0_resdetection_p_vsync)) begin
		soc_videooverlaysoc_hdmi_in0_resdetection_vcounter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in0_resdetection_pn_de) begin
			soc_videooverlaysoc_hdmi_in0_resdetection_vcounter <= (soc_videooverlaysoc_hdmi_in0_resdetection_vcounter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in0_resdetection_valid_i) begin
		if (soc_videooverlaysoc_hdmi_in0_resdetection_p_vsync) begin
			soc_videooverlaysoc_hdmi_in0_resdetection_vcounter_st <= soc_videooverlaysoc_hdmi_in0_resdetection_vcounter;
		end
	end else begin
		soc_videooverlaysoc_hdmi_in0_resdetection_vcounter_st <= 1'd0;
	end
	if (hdmi_in0_pix_rst) begin
		soc_videooverlaysoc_hdmi_in0_charsync0_synced <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_charsync0_data <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_charsync0_raw_data1 <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_charsync0_found_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_charsync0_control_counter <= 3'd0;
		soc_videooverlaysoc_hdmi_in0_charsync0_previous_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_charsync0_word_sel <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_data_r <= 9'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_transition_count <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_is_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_is_error <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_period_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_period_done <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_wer_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_r <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_r_updated <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding0_valid_o <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding0_output_raw <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_decoding0_output_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_decoding0_output_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_decoding0_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_charsync1_synced <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_charsync1_data <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_charsync1_raw_data1 <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_charsync1_found_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_charsync1_control_counter <= 3'd0;
		soc_videooverlaysoc_hdmi_in0_charsync1_previous_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_charsync1_word_sel <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_data_r <= 9'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_transition_count <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_is_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_is_error <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_period_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_period_done <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_wer_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_r <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_r_updated <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding1_valid_o <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding1_output_raw <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_decoding1_output_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_decoding1_output_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_decoding1_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_charsync2_synced <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_charsync2_data <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_charsync2_raw_data1 <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_charsync2_found_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_charsync2_control_counter <= 3'd0;
		soc_videooverlaysoc_hdmi_in0_charsync2_previous_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_charsync2_word_sel <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_data_r <= 9'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_transition_count <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_is_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_is_error <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_period_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_period_done <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_wer_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_r <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_r_updated <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding2_valid_o <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decoding2_output_raw <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_decoding2_output_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_decoding2_output_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_decoding2_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_chansync_chan_synced <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_produce <= 3'd0;
		soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_consume <= 3'd0;
		soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_produce <= 3'd0;
		soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_consume <= 3'd0;
		soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_produce <= 3'd0;
		soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_consume <= 3'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_de_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_syncpol_valid_o <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_syncpol_r <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_syncpol_g <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_syncpol_b <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_syncpol_de_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_syncpol_c_polarity <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_syncpol_c_out <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s0 <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s1 <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s2 <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_data0_timingdelay_next_s3 <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s0 <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s1 <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s2 <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_data1_timingdelay_next_s3 <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s0 <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s1 <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s2 <= 2'd0;
		soc_videooverlaysoc_hdmi_in0_data2_timingdelay_next_s3 <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_resdetection_de_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_resdetection_hcounter <= 11'd0;
		soc_videooverlaysoc_hdmi_in0_resdetection_hcounter_st <= 11'd0;
		soc_videooverlaysoc_hdmi_in0_resdetection_vsync_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_resdetection_vcounter <= 11'd0;
		soc_videooverlaysoc_hdmi_in0_resdetection_vcounter_st <= 11'd0;
		vns_clockdomainsrenamer0_state0 <= 3'd0;
	end
	vns_xilinxmultiregimpl37_regs0 <= soc_videooverlaysoc_hdmi_in0_decode_terc4_storage;
	vns_xilinxmultiregimpl37_regs1 <= vns_xilinxmultiregimpl37_regs0;
end

always @(posedge hdmi_in0_pix1p25x_clk) begin
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture0_reset_lateness) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_lateness <= 8'd128;
	end else begin
		if (((~soc_videooverlaysoc_hdmi_in0_s7datacapture0_too_late) & (~soc_videooverlaysoc_hdmi_in0_s7datacapture0_too_early))) begin
			if (soc_videooverlaysoc_hdmi_in0_s7datacapture0_dec) begin
				soc_videooverlaysoc_hdmi_in0_s7datacapture0_lateness <= (soc_videooverlaysoc_hdmi_in0_s7datacapture0_lateness + 1'd1);
			end
			if (soc_videooverlaysoc_hdmi_in0_s7datacapture0_inc) begin
				soc_videooverlaysoc_hdmi_in0_s7datacapture0_lateness <= (soc_videooverlaysoc_hdmi_in0_s7datacapture0_lateness - 1'd1);
			end
		end
	end
	soc_videooverlaysoc_hdmi_in0_s7datacapture0_mdata_d <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_mdata;
	soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_o;
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture1_reset_lateness) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_lateness <= 8'd128;
	end else begin
		if (((~soc_videooverlaysoc_hdmi_in0_s7datacapture1_too_late) & (~soc_videooverlaysoc_hdmi_in0_s7datacapture1_too_early))) begin
			if (soc_videooverlaysoc_hdmi_in0_s7datacapture1_dec) begin
				soc_videooverlaysoc_hdmi_in0_s7datacapture1_lateness <= (soc_videooverlaysoc_hdmi_in0_s7datacapture1_lateness + 1'd1);
			end
			if (soc_videooverlaysoc_hdmi_in0_s7datacapture1_inc) begin
				soc_videooverlaysoc_hdmi_in0_s7datacapture1_lateness <= (soc_videooverlaysoc_hdmi_in0_s7datacapture1_lateness - 1'd1);
			end
		end
	end
	soc_videooverlaysoc_hdmi_in0_s7datacapture1_mdata_d <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_mdata;
	soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_o;
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture2_reset_lateness) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_lateness <= 8'd128;
	end else begin
		if (((~soc_videooverlaysoc_hdmi_in0_s7datacapture2_too_late) & (~soc_videooverlaysoc_hdmi_in0_s7datacapture2_too_early))) begin
			if (soc_videooverlaysoc_hdmi_in0_s7datacapture2_dec) begin
				soc_videooverlaysoc_hdmi_in0_s7datacapture2_lateness <= (soc_videooverlaysoc_hdmi_in0_s7datacapture2_lateness + 1'd1);
			end
			if (soc_videooverlaysoc_hdmi_in0_s7datacapture2_inc) begin
				soc_videooverlaysoc_hdmi_in0_s7datacapture2_lateness <= (soc_videooverlaysoc_hdmi_in0_s7datacapture2_lateness - 1'd1);
			end
		end
	end
	soc_videooverlaysoc_hdmi_in0_s7datacapture2_mdata_d <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_mdata;
	soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_o;
	if (hdmi_in0_pix1p25x_rst) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_mdata_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_lateness <= 8'd128;
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_mdata_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_lateness <= 8'd128;
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_mdata_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_lateness <= 8'd128;
	end
	vns_xilinxmultiregimpl6_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_i;
	vns_xilinxmultiregimpl6_regs1 <= vns_xilinxmultiregimpl6_regs0;
	vns_xilinxmultiregimpl7_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_i;
	vns_xilinxmultiregimpl7_regs1 <= vns_xilinxmultiregimpl7_regs0;
	vns_xilinxmultiregimpl8_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_i;
	vns_xilinxmultiregimpl8_regs1 <= vns_xilinxmultiregimpl8_regs0;
	vns_xilinxmultiregimpl9_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_i;
	vns_xilinxmultiregimpl9_regs1 <= vns_xilinxmultiregimpl9_regs0;
	vns_xilinxmultiregimpl10_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_i;
	vns_xilinxmultiregimpl10_regs1 <= vns_xilinxmultiregimpl10_regs0;
	vns_xilinxmultiregimpl12_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_i;
	vns_xilinxmultiregimpl12_regs1 <= vns_xilinxmultiregimpl12_regs0;
	vns_xilinxmultiregimpl16_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_i;
	vns_xilinxmultiregimpl16_regs1 <= vns_xilinxmultiregimpl16_regs0;
	vns_xilinxmultiregimpl17_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_i;
	vns_xilinxmultiregimpl17_regs1 <= vns_xilinxmultiregimpl17_regs0;
	vns_xilinxmultiregimpl18_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_i;
	vns_xilinxmultiregimpl18_regs1 <= vns_xilinxmultiregimpl18_regs0;
	vns_xilinxmultiregimpl19_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_i;
	vns_xilinxmultiregimpl19_regs1 <= vns_xilinxmultiregimpl19_regs0;
	vns_xilinxmultiregimpl20_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_i;
	vns_xilinxmultiregimpl20_regs1 <= vns_xilinxmultiregimpl20_regs0;
	vns_xilinxmultiregimpl22_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_i;
	vns_xilinxmultiregimpl22_regs1 <= vns_xilinxmultiregimpl22_regs0;
	vns_xilinxmultiregimpl26_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_i;
	vns_xilinxmultiregimpl26_regs1 <= vns_xilinxmultiregimpl26_regs0;
	vns_xilinxmultiregimpl27_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_i;
	vns_xilinxmultiregimpl27_regs1 <= vns_xilinxmultiregimpl27_regs0;
	vns_xilinxmultiregimpl28_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_i;
	vns_xilinxmultiregimpl28_regs1 <= vns_xilinxmultiregimpl28_regs0;
	vns_xilinxmultiregimpl29_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_i;
	vns_xilinxmultiregimpl29_regs1 <= vns_xilinxmultiregimpl29_regs0;
	vns_xilinxmultiregimpl30_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_i;
	vns_xilinxmultiregimpl30_regs1 <= vns_xilinxmultiregimpl30_regs0;
	vns_xilinxmultiregimpl32_regs0 <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_i;
	vns_xilinxmultiregimpl32_regs1 <= vns_xilinxmultiregimpl32_regs0;
end

always @(posedge hdmi_in1_data0_cap_read_clk) begin
	soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst_read <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst;
	soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_rd <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr;
	if ((soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rdpointer == 3'd7)) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rdpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rdpointer <= (soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rdpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rdpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_rd[9:0];
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_rd[19:10];
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_rd[29:20];
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_rd[39:30];
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_rd[49:40];
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_rd[59:50];
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_rd[69:60];
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_rd[79:70];
		end
	endcase
	if (hdmi_in1_data0_cap_read_rst) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst_read <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge hdmi_in1_data0_cap_write_clk) begin
	soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst_write <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst;
	if ((soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_wrpointer == 4'd9)) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_wrpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_wrpointer <= (soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_wrpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_wrpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr[7:0] <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr[15:8] <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr[23:16] <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr[31:24] <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr[39:32] <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr[47:40] <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr[55:48] <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr[63:56] <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
		end
		4'd8: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr[71:64] <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
		end
		4'd9: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_storage_wr[79:72] <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_i;
		end
	endcase
	if (hdmi_in1_data0_cap_write_rst) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_rst_write <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge hdmi_in1_data1_cap_read_clk) begin
	soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst_read <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst;
	soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_rd <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr;
	if ((soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rdpointer == 3'd7)) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rdpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rdpointer <= (soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rdpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rdpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_rd[9:0];
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_rd[19:10];
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_rd[29:20];
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_rd[39:30];
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_rd[49:40];
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_rd[59:50];
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_rd[69:60];
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_rd[79:70];
		end
	endcase
	if (hdmi_in1_data1_cap_read_rst) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst_read <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge hdmi_in1_data1_cap_write_clk) begin
	soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst_write <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst;
	if ((soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_wrpointer == 4'd9)) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_wrpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_wrpointer <= (soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_wrpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_wrpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr[7:0] <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr[15:8] <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr[23:16] <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr[31:24] <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr[39:32] <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr[47:40] <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr[55:48] <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr[63:56] <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
		end
		4'd8: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr[71:64] <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
		end
		4'd9: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_storage_wr[79:72] <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_i;
		end
	endcase
	if (hdmi_in1_data1_cap_write_rst) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_rst_write <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge hdmi_in1_data2_cap_read_clk) begin
	soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst_read <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst;
	soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_rd <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr;
	if ((soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rdpointer == 3'd7)) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rdpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rdpointer <= (soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rdpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rdpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_rd[9:0];
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_rd[19:10];
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_rd[29:20];
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_rd[39:30];
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_rd[49:40];
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_rd[59:50];
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_rd[69:60];
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_o <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_rd[79:70];
		end
	endcase
	if (hdmi_in1_data2_cap_read_rst) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst_read <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge hdmi_in1_data2_cap_write_clk) begin
	soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst_write <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst;
	if ((soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_wrpointer == 4'd9)) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_wrpointer <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_wrpointer <= (soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_wrpointer + 1'd1);
	end
	case (soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_wrpointer)
		1'd0: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr[7:0] <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
		end
		1'd1: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr[15:8] <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
		end
		2'd2: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr[23:16] <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
		end
		2'd3: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr[31:24] <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
		end
		3'd4: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr[39:32] <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
		end
		3'd5: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr[47:40] <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
		end
		3'd6: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr[55:48] <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
		end
		3'd7: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr[63:56] <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
		end
		4'd8: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr[71:64] <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
		end
		4'd9: begin
			soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_storage_wr[79:72] <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_i;
		end
	endcase
	if (hdmi_in1_data2_cap_write_rst) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_rst_write <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge hdmi_in1_freq_fmeter_clk) begin
	soc_videooverlaysoc_hdmi_in1_freq_q_binary <= soc_videooverlaysoc_hdmi_in1_freq_q_next_binary;
	soc_videooverlaysoc_hdmi_in1_freq_q <= soc_videooverlaysoc_hdmi_in1_freq_q_next;
end

always @(posedge hdmi_in1_pix_clk) begin
	soc_videooverlaysoc_hdmi_in1_charsync0_raw_data1 <= soc_videooverlaysoc_hdmi_in1_charsync0_raw_data;
	soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd0;
	if (((((soc_videooverlaysoc_hdmi_in1_charsync0_raw[9:0] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[9:0] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[9:0] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[9:0] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 1'd0;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync0_raw[10:1] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[10:1] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[10:1] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[10:1] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 1'd1;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync0_raw[11:2] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[11:2] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[11:2] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[11:2] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 2'd2;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync0_raw[12:3] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[12:3] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[12:3] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[12:3] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 2'd3;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync0_raw[13:4] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[13:4] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[13:4] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[13:4] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 3'd4;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync0_raw[14:5] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[14:5] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[14:5] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[14:5] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 3'd5;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync0_raw[15:6] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[15:6] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[15:6] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[15:6] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 3'd6;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync0_raw[16:7] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[16:7] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[16:7] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[16:7] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 3'd7;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync0_raw[17:8] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[17:8] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[17:8] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[17:8] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 4'd8;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync0_raw[18:9] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[18:9] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[18:9] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync0_raw[18:9] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in1_charsync0_found_control & (soc_videooverlaysoc_hdmi_in1_charsync0_control_position == soc_videooverlaysoc_hdmi_in1_charsync0_previous_control_position))) begin
		if ((soc_videooverlaysoc_hdmi_in1_charsync0_control_counter == 3'd7)) begin
			soc_videooverlaysoc_hdmi_in1_charsync0_control_counter <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_charsync0_synced <= 1'd1;
			soc_videooverlaysoc_hdmi_in1_charsync0_word_sel <= soc_videooverlaysoc_hdmi_in1_charsync0_control_position;
		end else begin
			soc_videooverlaysoc_hdmi_in1_charsync0_control_counter <= (soc_videooverlaysoc_hdmi_in1_charsync0_control_counter + 1'd1);
		end
	end else begin
		soc_videooverlaysoc_hdmi_in1_charsync0_control_counter <= 1'd0;
	end
	soc_videooverlaysoc_hdmi_in1_charsync0_previous_control_position <= soc_videooverlaysoc_hdmi_in1_charsync0_control_position;
	soc_videooverlaysoc_hdmi_in1_charsync0_data <= (soc_videooverlaysoc_hdmi_in1_charsync0_raw >>> soc_videooverlaysoc_hdmi_in1_charsync0_word_sel);
	soc_videooverlaysoc_hdmi_in1_wer0_data_r <= soc_videooverlaysoc_hdmi_in1_wer0_data[8:0];
	soc_videooverlaysoc_hdmi_in1_wer0_transition_count <= (((((((soc_videooverlaysoc_hdmi_in1_wer0_transitions[0] + soc_videooverlaysoc_hdmi_in1_wer0_transitions[1]) + soc_videooverlaysoc_hdmi_in1_wer0_transitions[2]) + soc_videooverlaysoc_hdmi_in1_wer0_transitions[3]) + soc_videooverlaysoc_hdmi_in1_wer0_transitions[4]) + soc_videooverlaysoc_hdmi_in1_wer0_transitions[5]) + soc_videooverlaysoc_hdmi_in1_wer0_transitions[6]) + soc_videooverlaysoc_hdmi_in1_wer0_transitions[7]);
	soc_videooverlaysoc_hdmi_in1_wer0_is_control <= ((((soc_videooverlaysoc_hdmi_in1_wer0_data_r == 10'd852) | (soc_videooverlaysoc_hdmi_in1_wer0_data_r == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_wer0_data_r == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_wer0_data_r == 10'd683));
	soc_videooverlaysoc_hdmi_in1_wer0_is_error <= ((soc_videooverlaysoc_hdmi_in1_wer0_transition_count > 3'd4) & (~soc_videooverlaysoc_hdmi_in1_wer0_is_control));
	{soc_videooverlaysoc_hdmi_in1_wer0_period_done, soc_videooverlaysoc_hdmi_in1_wer0_period_counter} <= (soc_videooverlaysoc_hdmi_in1_wer0_period_counter + 1'd1);
	soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_r_updated <= soc_videooverlaysoc_hdmi_in1_wer0_period_done;
	if (soc_videooverlaysoc_hdmi_in1_wer0_period_done) begin
		soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_r <= soc_videooverlaysoc_hdmi_in1_wer0_wer_counter;
		soc_videooverlaysoc_hdmi_in1_wer0_wer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_wer0_is_error) begin
			soc_videooverlaysoc_hdmi_in1_wer0_wer_counter <= (soc_videooverlaysoc_hdmi_in1_wer0_wer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in1_wer0_i) begin
		soc_videooverlaysoc_hdmi_in1_wer0_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_wer0_toggle_i);
	end
	soc_videooverlaysoc_hdmi_in1_decoding0_output_de <= 1'd1;
	if ((soc_videooverlaysoc_hdmi_in1_decoding0_input == 10'd852)) begin
		soc_videooverlaysoc_hdmi_in1_decoding0_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding0_output_c <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decoding0_input == 8'd171)) begin
		soc_videooverlaysoc_hdmi_in1_decoding0_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding0_output_c <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decoding0_input == 9'd340)) begin
		soc_videooverlaysoc_hdmi_in1_decoding0_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding0_output_c <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decoding0_input == 10'd683)) begin
		soc_videooverlaysoc_hdmi_in1_decoding0_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding0_output_c <= 2'd3;
	end
	soc_videooverlaysoc_hdmi_in1_decoding0_output_raw <= soc_videooverlaysoc_hdmi_in1_decoding0_input;
	soc_videooverlaysoc_hdmi_in1_decoding0_output_d[0] <= (soc_videooverlaysoc_hdmi_in1_decoding0_input[0] ^ soc_videooverlaysoc_hdmi_in1_decoding0_input[9]);
	soc_videooverlaysoc_hdmi_in1_decoding0_output_d[1] <= ((soc_videooverlaysoc_hdmi_in1_decoding0_input[1] ^ soc_videooverlaysoc_hdmi_in1_decoding0_input[0]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding0_output_d[2] <= ((soc_videooverlaysoc_hdmi_in1_decoding0_input[2] ^ soc_videooverlaysoc_hdmi_in1_decoding0_input[1]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding0_output_d[3] <= ((soc_videooverlaysoc_hdmi_in1_decoding0_input[3] ^ soc_videooverlaysoc_hdmi_in1_decoding0_input[2]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding0_output_d[4] <= ((soc_videooverlaysoc_hdmi_in1_decoding0_input[4] ^ soc_videooverlaysoc_hdmi_in1_decoding0_input[3]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding0_output_d[5] <= ((soc_videooverlaysoc_hdmi_in1_decoding0_input[5] ^ soc_videooverlaysoc_hdmi_in1_decoding0_input[4]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding0_output_d[6] <= ((soc_videooverlaysoc_hdmi_in1_decoding0_input[6] ^ soc_videooverlaysoc_hdmi_in1_decoding0_input[5]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding0_output_d[7] <= ((soc_videooverlaysoc_hdmi_in1_decoding0_input[7] ^ soc_videooverlaysoc_hdmi_in1_decoding0_input[6]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding0_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding0_valid_o <= soc_videooverlaysoc_hdmi_in1_decoding0_valid_i;
	soc_videooverlaysoc_hdmi_in1_charsync1_raw_data1 <= soc_videooverlaysoc_hdmi_in1_charsync1_raw_data;
	soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd0;
	if (((((soc_videooverlaysoc_hdmi_in1_charsync1_raw[9:0] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[9:0] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[9:0] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[9:0] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 1'd0;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync1_raw[10:1] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[10:1] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[10:1] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[10:1] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 1'd1;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync1_raw[11:2] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[11:2] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[11:2] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[11:2] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 2'd2;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync1_raw[12:3] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[12:3] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[12:3] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[12:3] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 2'd3;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync1_raw[13:4] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[13:4] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[13:4] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[13:4] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 3'd4;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync1_raw[14:5] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[14:5] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[14:5] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[14:5] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 3'd5;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync1_raw[15:6] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[15:6] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[15:6] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[15:6] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 3'd6;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync1_raw[16:7] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[16:7] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[16:7] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[16:7] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 3'd7;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync1_raw[17:8] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[17:8] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[17:8] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[17:8] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 4'd8;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync1_raw[18:9] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[18:9] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[18:9] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync1_raw[18:9] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in1_charsync1_found_control & (soc_videooverlaysoc_hdmi_in1_charsync1_control_position == soc_videooverlaysoc_hdmi_in1_charsync1_previous_control_position))) begin
		if ((soc_videooverlaysoc_hdmi_in1_charsync1_control_counter == 3'd7)) begin
			soc_videooverlaysoc_hdmi_in1_charsync1_control_counter <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_charsync1_synced <= 1'd1;
			soc_videooverlaysoc_hdmi_in1_charsync1_word_sel <= soc_videooverlaysoc_hdmi_in1_charsync1_control_position;
		end else begin
			soc_videooverlaysoc_hdmi_in1_charsync1_control_counter <= (soc_videooverlaysoc_hdmi_in1_charsync1_control_counter + 1'd1);
		end
	end else begin
		soc_videooverlaysoc_hdmi_in1_charsync1_control_counter <= 1'd0;
	end
	soc_videooverlaysoc_hdmi_in1_charsync1_previous_control_position <= soc_videooverlaysoc_hdmi_in1_charsync1_control_position;
	soc_videooverlaysoc_hdmi_in1_charsync1_data <= (soc_videooverlaysoc_hdmi_in1_charsync1_raw >>> soc_videooverlaysoc_hdmi_in1_charsync1_word_sel);
	soc_videooverlaysoc_hdmi_in1_wer1_data_r <= soc_videooverlaysoc_hdmi_in1_wer1_data[8:0];
	soc_videooverlaysoc_hdmi_in1_wer1_transition_count <= (((((((soc_videooverlaysoc_hdmi_in1_wer1_transitions[0] + soc_videooverlaysoc_hdmi_in1_wer1_transitions[1]) + soc_videooverlaysoc_hdmi_in1_wer1_transitions[2]) + soc_videooverlaysoc_hdmi_in1_wer1_transitions[3]) + soc_videooverlaysoc_hdmi_in1_wer1_transitions[4]) + soc_videooverlaysoc_hdmi_in1_wer1_transitions[5]) + soc_videooverlaysoc_hdmi_in1_wer1_transitions[6]) + soc_videooverlaysoc_hdmi_in1_wer1_transitions[7]);
	soc_videooverlaysoc_hdmi_in1_wer1_is_control <= ((((soc_videooverlaysoc_hdmi_in1_wer1_data_r == 10'd852) | (soc_videooverlaysoc_hdmi_in1_wer1_data_r == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_wer1_data_r == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_wer1_data_r == 10'd683));
	soc_videooverlaysoc_hdmi_in1_wer1_is_error <= ((soc_videooverlaysoc_hdmi_in1_wer1_transition_count > 3'd4) & (~soc_videooverlaysoc_hdmi_in1_wer1_is_control));
	{soc_videooverlaysoc_hdmi_in1_wer1_period_done, soc_videooverlaysoc_hdmi_in1_wer1_period_counter} <= (soc_videooverlaysoc_hdmi_in1_wer1_period_counter + 1'd1);
	soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_r_updated <= soc_videooverlaysoc_hdmi_in1_wer1_period_done;
	if (soc_videooverlaysoc_hdmi_in1_wer1_period_done) begin
		soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_r <= soc_videooverlaysoc_hdmi_in1_wer1_wer_counter;
		soc_videooverlaysoc_hdmi_in1_wer1_wer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_wer1_is_error) begin
			soc_videooverlaysoc_hdmi_in1_wer1_wer_counter <= (soc_videooverlaysoc_hdmi_in1_wer1_wer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in1_wer1_i) begin
		soc_videooverlaysoc_hdmi_in1_wer1_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_wer1_toggle_i);
	end
	soc_videooverlaysoc_hdmi_in1_decoding1_output_de <= 1'd1;
	if ((soc_videooverlaysoc_hdmi_in1_decoding1_input == 10'd852)) begin
		soc_videooverlaysoc_hdmi_in1_decoding1_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding1_output_c <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decoding1_input == 8'd171)) begin
		soc_videooverlaysoc_hdmi_in1_decoding1_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding1_output_c <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decoding1_input == 9'd340)) begin
		soc_videooverlaysoc_hdmi_in1_decoding1_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding1_output_c <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decoding1_input == 10'd683)) begin
		soc_videooverlaysoc_hdmi_in1_decoding1_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding1_output_c <= 2'd3;
	end
	soc_videooverlaysoc_hdmi_in1_decoding1_output_raw <= soc_videooverlaysoc_hdmi_in1_decoding1_input;
	soc_videooverlaysoc_hdmi_in1_decoding1_output_d[0] <= (soc_videooverlaysoc_hdmi_in1_decoding1_input[0] ^ soc_videooverlaysoc_hdmi_in1_decoding1_input[9]);
	soc_videooverlaysoc_hdmi_in1_decoding1_output_d[1] <= ((soc_videooverlaysoc_hdmi_in1_decoding1_input[1] ^ soc_videooverlaysoc_hdmi_in1_decoding1_input[0]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding1_output_d[2] <= ((soc_videooverlaysoc_hdmi_in1_decoding1_input[2] ^ soc_videooverlaysoc_hdmi_in1_decoding1_input[1]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding1_output_d[3] <= ((soc_videooverlaysoc_hdmi_in1_decoding1_input[3] ^ soc_videooverlaysoc_hdmi_in1_decoding1_input[2]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding1_output_d[4] <= ((soc_videooverlaysoc_hdmi_in1_decoding1_input[4] ^ soc_videooverlaysoc_hdmi_in1_decoding1_input[3]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding1_output_d[5] <= ((soc_videooverlaysoc_hdmi_in1_decoding1_input[5] ^ soc_videooverlaysoc_hdmi_in1_decoding1_input[4]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding1_output_d[6] <= ((soc_videooverlaysoc_hdmi_in1_decoding1_input[6] ^ soc_videooverlaysoc_hdmi_in1_decoding1_input[5]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding1_output_d[7] <= ((soc_videooverlaysoc_hdmi_in1_decoding1_input[7] ^ soc_videooverlaysoc_hdmi_in1_decoding1_input[6]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding1_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding1_valid_o <= soc_videooverlaysoc_hdmi_in1_decoding1_valid_i;
	soc_videooverlaysoc_hdmi_in1_charsync2_raw_data1 <= soc_videooverlaysoc_hdmi_in1_charsync2_raw_data;
	soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd0;
	if (((((soc_videooverlaysoc_hdmi_in1_charsync2_raw[9:0] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[9:0] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[9:0] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[9:0] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 1'd0;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync2_raw[10:1] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[10:1] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[10:1] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[10:1] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 1'd1;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync2_raw[11:2] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[11:2] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[11:2] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[11:2] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 2'd2;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync2_raw[12:3] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[12:3] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[12:3] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[12:3] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 2'd3;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync2_raw[13:4] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[13:4] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[13:4] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[13:4] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 3'd4;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync2_raw[14:5] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[14:5] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[14:5] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[14:5] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 3'd5;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync2_raw[15:6] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[15:6] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[15:6] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[15:6] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 3'd6;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync2_raw[16:7] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[16:7] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[16:7] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[16:7] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 3'd7;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync2_raw[17:8] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[17:8] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[17:8] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[17:8] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 4'd8;
	end
	if (((((soc_videooverlaysoc_hdmi_in1_charsync2_raw[18:9] == 10'd852) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[18:9] == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[18:9] == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_charsync2_raw[18:9] == 10'd683))) begin
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in1_charsync2_found_control & (soc_videooverlaysoc_hdmi_in1_charsync2_control_position == soc_videooverlaysoc_hdmi_in1_charsync2_previous_control_position))) begin
		if ((soc_videooverlaysoc_hdmi_in1_charsync2_control_counter == 3'd7)) begin
			soc_videooverlaysoc_hdmi_in1_charsync2_control_counter <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_charsync2_synced <= 1'd1;
			soc_videooverlaysoc_hdmi_in1_charsync2_word_sel <= soc_videooverlaysoc_hdmi_in1_charsync2_control_position;
		end else begin
			soc_videooverlaysoc_hdmi_in1_charsync2_control_counter <= (soc_videooverlaysoc_hdmi_in1_charsync2_control_counter + 1'd1);
		end
	end else begin
		soc_videooverlaysoc_hdmi_in1_charsync2_control_counter <= 1'd0;
	end
	soc_videooverlaysoc_hdmi_in1_charsync2_previous_control_position <= soc_videooverlaysoc_hdmi_in1_charsync2_control_position;
	soc_videooverlaysoc_hdmi_in1_charsync2_data <= (soc_videooverlaysoc_hdmi_in1_charsync2_raw >>> soc_videooverlaysoc_hdmi_in1_charsync2_word_sel);
	soc_videooverlaysoc_hdmi_in1_wer2_data_r <= soc_videooverlaysoc_hdmi_in1_wer2_data[8:0];
	soc_videooverlaysoc_hdmi_in1_wer2_transition_count <= (((((((soc_videooverlaysoc_hdmi_in1_wer2_transitions[0] + soc_videooverlaysoc_hdmi_in1_wer2_transitions[1]) + soc_videooverlaysoc_hdmi_in1_wer2_transitions[2]) + soc_videooverlaysoc_hdmi_in1_wer2_transitions[3]) + soc_videooverlaysoc_hdmi_in1_wer2_transitions[4]) + soc_videooverlaysoc_hdmi_in1_wer2_transitions[5]) + soc_videooverlaysoc_hdmi_in1_wer2_transitions[6]) + soc_videooverlaysoc_hdmi_in1_wer2_transitions[7]);
	soc_videooverlaysoc_hdmi_in1_wer2_is_control <= ((((soc_videooverlaysoc_hdmi_in1_wer2_data_r == 10'd852) | (soc_videooverlaysoc_hdmi_in1_wer2_data_r == 8'd171)) | (soc_videooverlaysoc_hdmi_in1_wer2_data_r == 9'd340)) | (soc_videooverlaysoc_hdmi_in1_wer2_data_r == 10'd683));
	soc_videooverlaysoc_hdmi_in1_wer2_is_error <= ((soc_videooverlaysoc_hdmi_in1_wer2_transition_count > 3'd4) & (~soc_videooverlaysoc_hdmi_in1_wer2_is_control));
	{soc_videooverlaysoc_hdmi_in1_wer2_period_done, soc_videooverlaysoc_hdmi_in1_wer2_period_counter} <= (soc_videooverlaysoc_hdmi_in1_wer2_period_counter + 1'd1);
	soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_r_updated <= soc_videooverlaysoc_hdmi_in1_wer2_period_done;
	if (soc_videooverlaysoc_hdmi_in1_wer2_period_done) begin
		soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_r <= soc_videooverlaysoc_hdmi_in1_wer2_wer_counter;
		soc_videooverlaysoc_hdmi_in1_wer2_wer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_wer2_is_error) begin
			soc_videooverlaysoc_hdmi_in1_wer2_wer_counter <= (soc_videooverlaysoc_hdmi_in1_wer2_wer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in1_wer2_i) begin
		soc_videooverlaysoc_hdmi_in1_wer2_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_wer2_toggle_i);
	end
	soc_videooverlaysoc_hdmi_in1_decoding2_output_de <= 1'd1;
	if ((soc_videooverlaysoc_hdmi_in1_decoding2_input == 10'd852)) begin
		soc_videooverlaysoc_hdmi_in1_decoding2_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding2_output_c <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decoding2_input == 8'd171)) begin
		soc_videooverlaysoc_hdmi_in1_decoding2_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding2_output_c <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decoding2_input == 9'd340)) begin
		soc_videooverlaysoc_hdmi_in1_decoding2_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding2_output_c <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decoding2_input == 10'd683)) begin
		soc_videooverlaysoc_hdmi_in1_decoding2_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding2_output_c <= 2'd3;
	end
	soc_videooverlaysoc_hdmi_in1_decoding2_output_raw <= soc_videooverlaysoc_hdmi_in1_decoding2_input;
	soc_videooverlaysoc_hdmi_in1_decoding2_output_d[0] <= (soc_videooverlaysoc_hdmi_in1_decoding2_input[0] ^ soc_videooverlaysoc_hdmi_in1_decoding2_input[9]);
	soc_videooverlaysoc_hdmi_in1_decoding2_output_d[1] <= ((soc_videooverlaysoc_hdmi_in1_decoding2_input[1] ^ soc_videooverlaysoc_hdmi_in1_decoding2_input[0]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding2_output_d[2] <= ((soc_videooverlaysoc_hdmi_in1_decoding2_input[2] ^ soc_videooverlaysoc_hdmi_in1_decoding2_input[1]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding2_output_d[3] <= ((soc_videooverlaysoc_hdmi_in1_decoding2_input[3] ^ soc_videooverlaysoc_hdmi_in1_decoding2_input[2]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding2_output_d[4] <= ((soc_videooverlaysoc_hdmi_in1_decoding2_input[4] ^ soc_videooverlaysoc_hdmi_in1_decoding2_input[3]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding2_output_d[5] <= ((soc_videooverlaysoc_hdmi_in1_decoding2_input[5] ^ soc_videooverlaysoc_hdmi_in1_decoding2_input[4]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding2_output_d[6] <= ((soc_videooverlaysoc_hdmi_in1_decoding2_input[6] ^ soc_videooverlaysoc_hdmi_in1_decoding2_input[5]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding2_output_d[7] <= ((soc_videooverlaysoc_hdmi_in1_decoding2_input[7] ^ soc_videooverlaysoc_hdmi_in1_decoding2_input[6]) ^ (~soc_videooverlaysoc_hdmi_in1_decoding2_input[8]));
	soc_videooverlaysoc_hdmi_in1_decoding2_valid_o <= soc_videooverlaysoc_hdmi_in1_decoding2_valid_i;
	if ((~soc_videooverlaysoc_hdmi_in1_chansync_valid_i)) begin
		soc_videooverlaysoc_hdmi_in1_chansync_chan_synced <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_chansync_some_control) begin
			if (soc_videooverlaysoc_hdmi_in1_chansync_all_control) begin
				soc_videooverlaysoc_hdmi_in1_chansync_chan_synced <= 1'd1;
			end else begin
				soc_videooverlaysoc_hdmi_in1_chansync_chan_synced <= 1'd0;
			end
		end
	end
	soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_produce <= (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_produce + 1'd1);
	if (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_re) begin
		soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_consume <= (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_consume + 1'd1);
	end
	soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_produce <= (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_produce + 1'd1);
	if (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_re) begin
		soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_consume <= (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_consume + 1'd1);
	end
	soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_produce <= (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_produce + 1'd1);
	if (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_re) begin
		soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_consume <= (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_consume + 1'd1);
	end
	soc_videooverlaysoc_hdmi_in1_decode_terc4_de_r <= soc_videooverlaysoc_hdmi_in1_decode_terc4_data_in0_de;
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd668)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd611)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd740)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd738)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 2'd3;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 9'd369)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 3'd4;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 9'd286)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 3'd5;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 9'd398)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 3'd6;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 9'd316)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 3'd7;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd716)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd8;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 9'd313)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 9'd412)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd10;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd710)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd11;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd654)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd12;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd625)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd13;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 9'd355)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd14;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd707)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd15;
	end
	if (soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_valid_in) begin
		if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd852)) begin
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd1;
		end else begin
			if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 8'd171)) begin
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c <= 1'd1;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd1;
			end else begin
				if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 9'd340)) begin
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c <= 2'd2;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd1;
				end else begin
					if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd683)) begin
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c <= 2'd3;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd1;
					end else begin
						if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 9'd307)) begin
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c <= 1'd0;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd1;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd0;
						end else begin
							if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_data_in_raw == 10'd716)) begin
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd1;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd0;
							end else begin
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd1;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd0;
							end
						end
					end
				end
			end
		end
	end else begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd668)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd611)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd740)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd738)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 2'd3;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 9'd369)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 3'd4;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 9'd286)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 3'd5;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 9'd398)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 3'd6;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 9'd316)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 3'd7;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd716)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd8;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 9'd313)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 9'd412)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd10;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd710)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd11;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd654)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd12;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd625)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd13;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 9'd355)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd14;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd707)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd15;
	end
	if (soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_valid_in) begin
		if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd852)) begin
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd1;
		end else begin
			if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 8'd171)) begin
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c <= 1'd1;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd1;
			end else begin
				if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 9'd340)) begin
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c <= 2'd2;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd1;
				end else begin
					if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 10'd683)) begin
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c <= 2'd3;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd1;
					end else begin
						if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 9'd307)) begin
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c <= 1'd0;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd1;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd1;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd0;
						end else begin
							if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_data_in_raw == 9'd307)) begin
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd1;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd1;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd0;
							end else begin
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd1;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd0;
							end
						end
					end
				end
			end
		end
	end else begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd668)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 1'd0;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd611)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 1'd1;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd740)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 2'd2;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd738)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 2'd3;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 9'd369)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 3'd4;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 9'd286)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 3'd5;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 9'd398)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 3'd6;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 9'd316)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 3'd7;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd716)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd8;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 9'd313)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd9;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 9'd412)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd10;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd710)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd11;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd654)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd12;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd625)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd13;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 9'd355)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd14;
	end
	if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd707)) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd15;
	end
	if (soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_valid_in) begin
		if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd852)) begin
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
			soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd1;
		end else begin
			if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 8'd171)) begin
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c <= 1'd1;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
				soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd1;
			end else begin
				if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 9'd340)) begin
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c <= 2'd2;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
					soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd1;
				end else begin
					if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd683)) begin
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c <= 2'd3;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
						soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd1;
					end else begin
						if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 9'd307)) begin
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c <= 1'd0;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd1;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
							soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd0;
						end else begin
							if ((soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_data_in_raw == 10'd716)) begin
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd1;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd0;
							end else begin
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd1;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
								soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd0;
							end
						end
					end
				end
			end
		end
	end else begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd0;
	end
	vns_clockdomainsrenamer1_state0 <= vns_clockdomainsrenamer1_next_state0;
	soc_videooverlaysoc_hdmi_in1_syncpol_valid_o <= soc_videooverlaysoc_hdmi_in1_syncpol_valid_i;
	soc_videooverlaysoc_hdmi_in1_syncpol_r <= soc_videooverlaysoc_hdmi_in1_syncpol_data_in2_d;
	soc_videooverlaysoc_hdmi_in1_syncpol_g <= soc_videooverlaysoc_hdmi_in1_syncpol_data_in1_d;
	soc_videooverlaysoc_hdmi_in1_syncpol_b <= soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_d;
	soc_videooverlaysoc_hdmi_in1_syncpol_de_r <= soc_videooverlaysoc_hdmi_in1_syncpol_de_int;
	if (soc_videooverlaysoc_hdmi_in1_syncpol_de_rising) begin
		soc_videooverlaysoc_hdmi_in1_syncpol_c_polarity <= soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_c;
		soc_videooverlaysoc_hdmi_in1_syncpol_c_out <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in1_syncpol_c_out <= (soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_c ^ soc_videooverlaysoc_hdmi_in1_syncpol_c_polarity);
	end
	soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s0 <= soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_raw;
	soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s1 <= soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_d;
	soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s2 <= soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_c;
	soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s3 <= soc_videooverlaysoc_hdmi_in1_data0_timingdelay_sink_de;
	soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s0 <= soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_raw;
	soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s1 <= soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_d;
	soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s2 <= soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_c;
	soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s3 <= soc_videooverlaysoc_hdmi_in1_data1_timingdelay_sink_de;
	soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s0 <= soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_raw;
	soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s1 <= soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_d;
	soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s2 <= soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_c;
	soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s3 <= soc_videooverlaysoc_hdmi_in1_data2_timingdelay_sink_de;
	soc_videooverlaysoc_hdmi_in1_resdetection_de_r <= soc_videooverlaysoc_hdmi_in1_resdetection_de;
	if ((soc_videooverlaysoc_hdmi_in1_resdetection_valid_i & soc_videooverlaysoc_hdmi_in1_resdetection_de)) begin
		soc_videooverlaysoc_hdmi_in1_resdetection_hcounter <= (soc_videooverlaysoc_hdmi_in1_resdetection_hcounter + 1'd1);
	end else begin
		soc_videooverlaysoc_hdmi_in1_resdetection_hcounter <= 1'd0;
	end
	if (soc_videooverlaysoc_hdmi_in1_resdetection_valid_i) begin
		if (soc_videooverlaysoc_hdmi_in1_resdetection_pn_de) begin
			soc_videooverlaysoc_hdmi_in1_resdetection_hcounter_st <= soc_videooverlaysoc_hdmi_in1_resdetection_hcounter;
		end
	end else begin
		soc_videooverlaysoc_hdmi_in1_resdetection_hcounter_st <= 1'd0;
	end
	soc_videooverlaysoc_hdmi_in1_resdetection_vsync_r <= soc_videooverlaysoc_hdmi_in1_resdetection_vsync;
	if ((soc_videooverlaysoc_hdmi_in1_resdetection_valid_i & soc_videooverlaysoc_hdmi_in1_resdetection_p_vsync)) begin
		soc_videooverlaysoc_hdmi_in1_resdetection_vcounter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_resdetection_pn_de) begin
			soc_videooverlaysoc_hdmi_in1_resdetection_vcounter <= (soc_videooverlaysoc_hdmi_in1_resdetection_vcounter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in1_resdetection_valid_i) begin
		if (soc_videooverlaysoc_hdmi_in1_resdetection_p_vsync) begin
			soc_videooverlaysoc_hdmi_in1_resdetection_vcounter_st <= soc_videooverlaysoc_hdmi_in1_resdetection_vcounter;
		end
	end else begin
		soc_videooverlaysoc_hdmi_in1_resdetection_vcounter_st <= 1'd0;
	end
	soc_videooverlaysoc_hdmi_in1_frame_vsync_r <= soc_videooverlaysoc_hdmi_in1_frame_vsync;
	soc_videooverlaysoc_hdmi_in1_frame_cur_word_valid <= 1'd0;
	if (soc_videooverlaysoc_hdmi_in1_frame_new_frame) begin
		soc_videooverlaysoc_hdmi_in1_frame_cur_word_valid <= (soc_videooverlaysoc_hdmi_in1_frame_pack_counter == 3'd7);
		soc_videooverlaysoc_hdmi_in1_frame_pack_counter <= 1'd0;
	end else begin
		if ((soc_videooverlaysoc_hdmi_in1_frame_valid_i & soc_videooverlaysoc_hdmi_in1_frame_de)) begin
			if ((soc_videooverlaysoc_hdmi_in1_frame_pack_counter == 3'd7)) begin
				soc_videooverlaysoc_hdmi_in1_frame_cur_word[31:0] <= soc_videooverlaysoc_hdmi_in1_frame_encoded_pixel;
			end
			if ((soc_videooverlaysoc_hdmi_in1_frame_pack_counter == 3'd6)) begin
				soc_videooverlaysoc_hdmi_in1_frame_cur_word[63:32] <= soc_videooverlaysoc_hdmi_in1_frame_encoded_pixel;
			end
			if ((soc_videooverlaysoc_hdmi_in1_frame_pack_counter == 3'd5)) begin
				soc_videooverlaysoc_hdmi_in1_frame_cur_word[95:64] <= soc_videooverlaysoc_hdmi_in1_frame_encoded_pixel;
			end
			if ((soc_videooverlaysoc_hdmi_in1_frame_pack_counter == 3'd4)) begin
				soc_videooverlaysoc_hdmi_in1_frame_cur_word[127:96] <= soc_videooverlaysoc_hdmi_in1_frame_encoded_pixel;
			end
			if ((soc_videooverlaysoc_hdmi_in1_frame_pack_counter == 2'd3)) begin
				soc_videooverlaysoc_hdmi_in1_frame_cur_word[159:128] <= soc_videooverlaysoc_hdmi_in1_frame_encoded_pixel;
			end
			if ((soc_videooverlaysoc_hdmi_in1_frame_pack_counter == 2'd2)) begin
				soc_videooverlaysoc_hdmi_in1_frame_cur_word[191:160] <= soc_videooverlaysoc_hdmi_in1_frame_encoded_pixel;
			end
			if ((soc_videooverlaysoc_hdmi_in1_frame_pack_counter == 1'd1)) begin
				soc_videooverlaysoc_hdmi_in1_frame_cur_word[223:192] <= soc_videooverlaysoc_hdmi_in1_frame_encoded_pixel;
			end
			if ((soc_videooverlaysoc_hdmi_in1_frame_pack_counter == 1'd0)) begin
				soc_videooverlaysoc_hdmi_in1_frame_cur_word[255:224] <= soc_videooverlaysoc_hdmi_in1_frame_encoded_pixel;
			end
			soc_videooverlaysoc_hdmi_in1_frame_cur_word_valid <= (soc_videooverlaysoc_hdmi_in1_frame_pack_counter == 3'd7);
			soc_videooverlaysoc_hdmi_in1_frame_pack_counter <= (soc_videooverlaysoc_hdmi_in1_frame_pack_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in1_frame_new_frame) begin
		soc_videooverlaysoc_hdmi_in1_frame_sink_payload_sof <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_frame_cur_word_valid) begin
			soc_videooverlaysoc_hdmi_in1_frame_sink_payload_sof <= 1'd0;
		end
	end
	if ((soc_videooverlaysoc_hdmi_in1_frame_sink_valid & (~soc_videooverlaysoc_hdmi_in1_frame_sink_ready))) begin
		soc_videooverlaysoc_hdmi_in1_frame_pix_overflow <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_frame_pix_overflow_reset) begin
			soc_videooverlaysoc_hdmi_in1_frame_pix_overflow <= 1'd0;
		end
	end
	soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_binary <= soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_next_binary;
	soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q <= soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_next;
	soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_o;
	if (soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_i) begin
		soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_i);
	end
	if (hdmi_in1_pix_rst) begin
		soc_videooverlaysoc_hdmi_in1_charsync0_synced <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_charsync0_data <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_charsync0_raw_data1 <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_charsync0_found_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_charsync0_control_counter <= 3'd0;
		soc_videooverlaysoc_hdmi_in1_charsync0_previous_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_charsync0_word_sel <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_data_r <= 9'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_transition_count <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_is_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_is_error <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_period_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_period_done <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_wer_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_r <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_r_updated <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding0_valid_o <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding0_output_raw <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_decoding0_output_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_decoding0_output_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_decoding0_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_charsync1_synced <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_charsync1_data <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_charsync1_raw_data1 <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_charsync1_found_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_charsync1_control_counter <= 3'd0;
		soc_videooverlaysoc_hdmi_in1_charsync1_previous_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_charsync1_word_sel <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_data_r <= 9'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_transition_count <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_is_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_is_error <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_period_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_period_done <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_wer_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_r <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_r_updated <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding1_valid_o <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding1_output_raw <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_decoding1_output_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_decoding1_output_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_decoding1_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_charsync2_synced <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_charsync2_data <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_charsync2_raw_data1 <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_charsync2_found_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_charsync2_control_counter <= 3'd0;
		soc_videooverlaysoc_hdmi_in1_charsync2_previous_control_position <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_charsync2_word_sel <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_data_r <= 9'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_transition_count <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_is_control <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_is_error <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_period_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_period_done <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_wer_counter <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_r <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_r_updated <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding2_valid_o <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decoding2_output_raw <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_decoding2_output_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_decoding2_output_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_decoding2_output_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_chansync_chan_synced <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_produce <= 3'd0;
		soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_consume <= 3'd0;
		soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_produce <= 3'd0;
		soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_consume <= 3'd0;
		soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_produce <= 3'd0;
		soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_consume <= 3'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_de_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_c_valid <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel0_decval_payload_d <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_c_valid <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel1_decval_payload_d <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_dgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_vgb <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_c_valid <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_decodeterc4channel2_decval_payload_d <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_syncpol_valid_o <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_syncpol_r <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_syncpol_g <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_syncpol_b <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_syncpol_de_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_syncpol_c_polarity <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_syncpol_c_out <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s0 <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s1 <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s2 <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_data0_timingdelay_next_s3 <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s0 <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s1 <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s2 <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_data1_timingdelay_next_s3 <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s0 <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s1 <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s2 <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_data2_timingdelay_next_s3 <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_resdetection_de_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_resdetection_hcounter <= 11'd0;
		soc_videooverlaysoc_hdmi_in1_resdetection_hcounter_st <= 11'd0;
		soc_videooverlaysoc_hdmi_in1_resdetection_vsync_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_resdetection_vcounter <= 11'd0;
		soc_videooverlaysoc_hdmi_in1_resdetection_vcounter_st <= 11'd0;
		soc_videooverlaysoc_hdmi_in1_frame_vsync_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_frame_cur_word <= 256'd0;
		soc_videooverlaysoc_hdmi_in1_frame_cur_word_valid <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_frame_pack_counter <= 3'd0;
		soc_videooverlaysoc_hdmi_in1_frame_sink_payload_sof <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q <= 11'd0;
		soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q_binary <= 11'd0;
		soc_videooverlaysoc_hdmi_in1_frame_pix_overflow <= 1'd0;
		vns_clockdomainsrenamer1_state0 <= 3'd0;
	end
	vns_xilinxmultiregimpl75_regs0 <= soc_videooverlaysoc_hdmi_in1_decode_terc4_storage;
	vns_xilinxmultiregimpl75_regs1 <= vns_xilinxmultiregimpl75_regs0;
	vns_xilinxmultiregimpl79_regs0 <= soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q;
	vns_xilinxmultiregimpl79_regs1 <= vns_xilinxmultiregimpl79_regs0;
	vns_xilinxmultiregimpl81_regs0 <= soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_i;
	vns_xilinxmultiregimpl81_regs1 <= vns_xilinxmultiregimpl81_regs0;
end

always @(posedge hdmi_in1_pix1p25x_clk) begin
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture0_reset_lateness) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_lateness <= 8'd128;
	end else begin
		if (((~soc_videooverlaysoc_hdmi_in1_s7datacapture0_too_late) & (~soc_videooverlaysoc_hdmi_in1_s7datacapture0_too_early))) begin
			if (soc_videooverlaysoc_hdmi_in1_s7datacapture0_dec) begin
				soc_videooverlaysoc_hdmi_in1_s7datacapture0_lateness <= (soc_videooverlaysoc_hdmi_in1_s7datacapture0_lateness + 1'd1);
			end
			if (soc_videooverlaysoc_hdmi_in1_s7datacapture0_inc) begin
				soc_videooverlaysoc_hdmi_in1_s7datacapture0_lateness <= (soc_videooverlaysoc_hdmi_in1_s7datacapture0_lateness - 1'd1);
			end
		end
	end
	soc_videooverlaysoc_hdmi_in1_s7datacapture0_mdata_d <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_mdata;
	soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_o;
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture1_reset_lateness) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_lateness <= 8'd128;
	end else begin
		if (((~soc_videooverlaysoc_hdmi_in1_s7datacapture1_too_late) & (~soc_videooverlaysoc_hdmi_in1_s7datacapture1_too_early))) begin
			if (soc_videooverlaysoc_hdmi_in1_s7datacapture1_dec) begin
				soc_videooverlaysoc_hdmi_in1_s7datacapture1_lateness <= (soc_videooverlaysoc_hdmi_in1_s7datacapture1_lateness + 1'd1);
			end
			if (soc_videooverlaysoc_hdmi_in1_s7datacapture1_inc) begin
				soc_videooverlaysoc_hdmi_in1_s7datacapture1_lateness <= (soc_videooverlaysoc_hdmi_in1_s7datacapture1_lateness - 1'd1);
			end
		end
	end
	soc_videooverlaysoc_hdmi_in1_s7datacapture1_mdata_d <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_mdata;
	soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_o;
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture2_reset_lateness) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_lateness <= 8'd128;
	end else begin
		if (((~soc_videooverlaysoc_hdmi_in1_s7datacapture2_too_late) & (~soc_videooverlaysoc_hdmi_in1_s7datacapture2_too_early))) begin
			if (soc_videooverlaysoc_hdmi_in1_s7datacapture2_dec) begin
				soc_videooverlaysoc_hdmi_in1_s7datacapture2_lateness <= (soc_videooverlaysoc_hdmi_in1_s7datacapture2_lateness + 1'd1);
			end
			if (soc_videooverlaysoc_hdmi_in1_s7datacapture2_inc) begin
				soc_videooverlaysoc_hdmi_in1_s7datacapture2_lateness <= (soc_videooverlaysoc_hdmi_in1_s7datacapture2_lateness - 1'd1);
			end
		end
	end
	soc_videooverlaysoc_hdmi_in1_s7datacapture2_mdata_d <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_mdata;
	soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_o;
	soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_o;
	if (hdmi_in1_pix1p25x_rst) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_mdata_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_lateness <= 8'd128;
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_mdata_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_lateness <= 8'd128;
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_mdata_d <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_lateness <= 8'd128;
	end
	vns_xilinxmultiregimpl44_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_i;
	vns_xilinxmultiregimpl44_regs1 <= vns_xilinxmultiregimpl44_regs0;
	vns_xilinxmultiregimpl45_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_i;
	vns_xilinxmultiregimpl45_regs1 <= vns_xilinxmultiregimpl45_regs0;
	vns_xilinxmultiregimpl46_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_i;
	vns_xilinxmultiregimpl46_regs1 <= vns_xilinxmultiregimpl46_regs0;
	vns_xilinxmultiregimpl47_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_i;
	vns_xilinxmultiregimpl47_regs1 <= vns_xilinxmultiregimpl47_regs0;
	vns_xilinxmultiregimpl48_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_i;
	vns_xilinxmultiregimpl48_regs1 <= vns_xilinxmultiregimpl48_regs0;
	vns_xilinxmultiregimpl50_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_i;
	vns_xilinxmultiregimpl50_regs1 <= vns_xilinxmultiregimpl50_regs0;
	vns_xilinxmultiregimpl54_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_i;
	vns_xilinxmultiregimpl54_regs1 <= vns_xilinxmultiregimpl54_regs0;
	vns_xilinxmultiregimpl55_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_i;
	vns_xilinxmultiregimpl55_regs1 <= vns_xilinxmultiregimpl55_regs0;
	vns_xilinxmultiregimpl56_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_i;
	vns_xilinxmultiregimpl56_regs1 <= vns_xilinxmultiregimpl56_regs0;
	vns_xilinxmultiregimpl57_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_i;
	vns_xilinxmultiregimpl57_regs1 <= vns_xilinxmultiregimpl57_regs0;
	vns_xilinxmultiregimpl58_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_i;
	vns_xilinxmultiregimpl58_regs1 <= vns_xilinxmultiregimpl58_regs0;
	vns_xilinxmultiregimpl60_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_i;
	vns_xilinxmultiregimpl60_regs1 <= vns_xilinxmultiregimpl60_regs0;
	vns_xilinxmultiregimpl64_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_i;
	vns_xilinxmultiregimpl64_regs1 <= vns_xilinxmultiregimpl64_regs0;
	vns_xilinxmultiregimpl65_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_i;
	vns_xilinxmultiregimpl65_regs1 <= vns_xilinxmultiregimpl65_regs0;
	vns_xilinxmultiregimpl66_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_i;
	vns_xilinxmultiregimpl66_regs1 <= vns_xilinxmultiregimpl66_regs0;
	vns_xilinxmultiregimpl67_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_i;
	vns_xilinxmultiregimpl67_regs1 <= vns_xilinxmultiregimpl67_regs0;
	vns_xilinxmultiregimpl68_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_i;
	vns_xilinxmultiregimpl68_regs1 <= vns_xilinxmultiregimpl68_regs0;
	vns_xilinxmultiregimpl70_regs0 <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_i;
	vns_xilinxmultiregimpl70_regs1 <= vns_xilinxmultiregimpl70_regs0;
end

always @(posedge pix_o_clk) begin
	soc_videooverlaysoc_hdmi_in0_timing_payload_de <= soc_videooverlaysoc_hdmi_in0_syncpol_de;
	soc_videooverlaysoc_hdmi_in0_timing_payload_hsync <= soc_videooverlaysoc_hdmi_in0_syncpol_hsync;
	soc_videooverlaysoc_hdmi_in0_timing_payload_vsync <= soc_videooverlaysoc_hdmi_in0_syncpol_vsync;
	if (soc_videooverlaysoc_hdmi_in0_syncpol_valid_o) begin
		soc_videooverlaysoc_hdmi_in0_timing_valid <= 1'd1;
	end else begin
		soc_videooverlaysoc_hdmi_in0_timing_valid <= 1'd0;
	end
	soc_videooverlaysoc_core_source_valid_d <= soc_videooverlaysoc_hdmi_core_out0_source_source_valid;
	soc_videooverlaysoc_core_source_data_d <= soc_videooverlaysoc_hdmi_core_out0_source_source_payload_data;
	soc_videooverlaysoc_Aksv14_r <= soc_videooverlaysoc_Aksv14;
	soc_videooverlaysoc_hdcp_Aksv14_write <= (soc_videooverlaysoc_Aksv14 & (~soc_videooverlaysoc_Aksv14_r));
	soc_videooverlaysoc_hdcp_hdcp_ena <= (soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_video | soc_videooverlaysoc_hdmi_in0_decode_terc4_encrypting_data);
	soc_videooverlaysoc_hdcp_hpd <= hdmi_in0_hpd_notif;
	soc_videooverlaysoc_hdcp_An <= soc_videooverlaysoc_i2c_snoop_An;
	soc_videooverlaysoc_hdcp_ctl_code <= soc_videooverlaysoc_hdmi_in0_decode_terc4_ctl_code;
	soc_videooverlaysoc_c0_next0 <= soc_videooverlaysoc_c0;
	soc_videooverlaysoc_c1_next0 <= soc_videooverlaysoc_c1;
	soc_videooverlaysoc_c2_next0 <= soc_videooverlaysoc_c2;
	soc_videooverlaysoc_c0_next1 <= soc_videooverlaysoc_c0_next0;
	soc_videooverlaysoc_c1_next1 <= soc_videooverlaysoc_c1_next0;
	soc_videooverlaysoc_c2_next1 <= soc_videooverlaysoc_c2_next0;
	soc_videooverlaysoc_c0_next2 <= soc_videooverlaysoc_c0_next1;
	soc_videooverlaysoc_c1_next2 <= soc_videooverlaysoc_c1_next1;
	soc_videooverlaysoc_c2_next2 <= soc_videooverlaysoc_c2_next1;
	soc_videooverlaysoc_c0_next3 <= soc_videooverlaysoc_c0_next2;
	soc_videooverlaysoc_c1_next3 <= soc_videooverlaysoc_c1_next2;
	soc_videooverlaysoc_c2_next3 <= soc_videooverlaysoc_c2_next2;
	soc_videooverlaysoc_c0_next4 <= soc_videooverlaysoc_c0_next3;
	soc_videooverlaysoc_c1_next4 <= soc_videooverlaysoc_c1_next3;
	soc_videooverlaysoc_c2_next4 <= soc_videooverlaysoc_c2_next3;
	soc_videooverlaysoc_c0_next5 <= soc_videooverlaysoc_c0_next4;
	soc_videooverlaysoc_c1_next5 <= soc_videooverlaysoc_c1_next4;
	soc_videooverlaysoc_c2_next5 <= soc_videooverlaysoc_c2_next4;
	soc_videooverlaysoc_c0_pix_o <= soc_videooverlaysoc_c0_next5;
	soc_videooverlaysoc_c1_pix_o <= soc_videooverlaysoc_c1_next5;
	soc_videooverlaysoc_c2_pix_o <= soc_videooverlaysoc_c2_next5;
	if ((((soc_videooverlaysoc_rect_on0 & (soc_videooverlaysoc_hdmi_out0_rgb_d_payload_r >= soc_videooverlaysoc_rect_thresh)) & (soc_videooverlaysoc_hdmi_out0_rgb_d_payload_g >= soc_videooverlaysoc_rect_thresh)) & (soc_videooverlaysoc_hdmi_out0_rgb_d_payload_b >= soc_videooverlaysoc_rect_thresh))) begin
		soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c0 <= soc_videooverlaysoc_encoder2_out;
		soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c1 <= soc_videooverlaysoc_encoder1_out;
		soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c2 <= soc_videooverlaysoc_encoder0_out;
	end else begin
		soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c0 <= soc_videooverlaysoc_c0_pix_o;
		soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c1 <= soc_videooverlaysoc_c1_pix_o;
		soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c2 <= soc_videooverlaysoc_c2_pix_o;
	end
	soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_binary <= soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_next_binary;
	soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q <= soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_next;
	soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_binary <= soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next_binary;
	soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q <= soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_next;
	if (soc_videooverlaysoc_out_dram_port_counter_ce) begin
		soc_videooverlaysoc_out_dram_port_counter <= (soc_videooverlaysoc_out_dram_port_counter + 1'd1);
	end
	if ((soc_videooverlaysoc_out_dram_port_rdata_converter_source_valid & soc_videooverlaysoc_out_dram_port_rdata_converter_source_ready)) begin
		soc_videooverlaysoc_out_dram_port_rdata_chunk <= {soc_videooverlaysoc_out_dram_port_rdata_chunk[6:0], soc_videooverlaysoc_out_dram_port_rdata_chunk[7]};
	end
	if (((soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_we & soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_writable) & (~soc_videooverlaysoc_out_dram_port_cmd_buffer_replace))) begin
		soc_videooverlaysoc_out_dram_port_cmd_buffer_produce <= (soc_videooverlaysoc_out_dram_port_cmd_buffer_produce + 1'd1);
	end
	if (soc_videooverlaysoc_out_dram_port_cmd_buffer_do_read) begin
		soc_videooverlaysoc_out_dram_port_cmd_buffer_consume <= (soc_videooverlaysoc_out_dram_port_cmd_buffer_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_we & soc_videooverlaysoc_out_dram_port_cmd_buffer_syncfifo_writable) & (~soc_videooverlaysoc_out_dram_port_cmd_buffer_replace))) begin
		if ((~soc_videooverlaysoc_out_dram_port_cmd_buffer_do_read)) begin
			soc_videooverlaysoc_out_dram_port_cmd_buffer_level <= (soc_videooverlaysoc_out_dram_port_cmd_buffer_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_out_dram_port_cmd_buffer_do_read) begin
			soc_videooverlaysoc_out_dram_port_cmd_buffer_level <= (soc_videooverlaysoc_out_dram_port_cmd_buffer_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_out_dram_port_rdata_buffer_pipe_ce) begin
		soc_videooverlaysoc_out_dram_port_rdata_buffer_valid_n <= soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_valid;
	end
	if (soc_videooverlaysoc_out_dram_port_rdata_buffer_pipe_ce) begin
		soc_videooverlaysoc_out_dram_port_rdata_buffer_first_n <= (soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_valid & soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_first);
		soc_videooverlaysoc_out_dram_port_rdata_buffer_last_n <= (soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_valid & soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_last);
	end
	if (soc_videooverlaysoc_out_dram_port_rdata_buffer_pipe_ce) begin
		soc_videooverlaysoc_out_dram_port_rdata_buffer_source_payload_data <= soc_videooverlaysoc_out_dram_port_rdata_buffer_sink_payload_data;
	end
	if ((soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_valid & soc_videooverlaysoc_out_dram_port_rdata_converter_converter_source_ready)) begin
		if (soc_videooverlaysoc_out_dram_port_rdata_converter_converter_last) begin
			soc_videooverlaysoc_out_dram_port_rdata_converter_converter_mux <= 1'd0;
		end else begin
			soc_videooverlaysoc_out_dram_port_rdata_converter_converter_mux <= (soc_videooverlaysoc_out_dram_port_rdata_converter_converter_mux + 1'd1);
		end
	end
	soc_videooverlaysoc_hdmi_in0_syncpol_c0 <= soc_videooverlaysoc_hdmi_in0_syncpol_data_in0_raw;
	soc_videooverlaysoc_hdmi_in0_syncpol_c1 <= soc_videooverlaysoc_hdmi_in0_syncpol_data_in1_raw;
	soc_videooverlaysoc_hdmi_in0_syncpol_c2 <= soc_videooverlaysoc_hdmi_in0_syncpol_data_in2_raw;
	soc_videooverlaysoc_hdmi_out0_clk_gen_ce <= (~pix_o_rst);
	soc_videooverlaysoc_hdmi_out0_phy_es0_ce <= (~pix_o_rst);
	soc_videooverlaysoc_hdmi_out0_phy_es1_ce <= (~pix_o_rst);
	soc_videooverlaysoc_hdmi_out0_phy_es2_ce <= (~pix_o_rst);
	soc_videooverlaysoc_hdmi_in1_syncpol_c0 <= soc_videooverlaysoc_hdmi_in1_syncpol_data_in0_raw;
	soc_videooverlaysoc_hdmi_in1_syncpol_c1 <= soc_videooverlaysoc_hdmi_in1_syncpol_data_in1_raw;
	soc_videooverlaysoc_hdmi_in1_syncpol_c2 <= soc_videooverlaysoc_hdmi_in1_syncpol_data_in2_raw;
	if (soc_videooverlaysoc_hdmi_core_out0_underflow_enable) begin
		if ((~soc_videooverlaysoc_hdmi_core_out0_source_source_valid)) begin
			soc_videooverlaysoc_hdmi_core_out0_underflow_counter <= (soc_videooverlaysoc_hdmi_core_out0_underflow_counter + 1'd1);
		end
	end else begin
		soc_videooverlaysoc_hdmi_core_out0_underflow_counter <= 1'd0;
	end
	if (soc_videooverlaysoc_hdmi_core_out0_underflow_update) begin
		soc_videooverlaysoc_hdmi_core_out0_underflow_counter_status <= soc_videooverlaysoc_hdmi_core_out0_underflow_counter;
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_binary <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next_binary;
	soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_next;
	soc_videooverlaysoc_hdmi_core_out0_dmareader_v <= soc_videooverlaysoc_hdmi_in0_timing_payload_vsync;
	soc_videooverlaysoc_hdmi_core_out0_dmareader_v_r <= soc_videooverlaysoc_hdmi_core_out0_dmareader_v;
	soc_videooverlaysoc_hdmi_core_out0_dmareader_sof <= (soc_videooverlaysoc_hdmi_core_out0_dmareader_v & (~soc_videooverlaysoc_hdmi_core_out0_dmareader_v_r));
	if (soc_videooverlaysoc_hdmi_core_out0_dmareader_request_issued) begin
		if ((~soc_videooverlaysoc_hdmi_core_out0_dmareader_data_dequeued)) begin
			soc_videooverlaysoc_hdmi_core_out0_dmareader_rsv_level <= (soc_videooverlaysoc_hdmi_core_out0_dmareader_rsv_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_hdmi_core_out0_dmareader_data_dequeued) begin
			soc_videooverlaysoc_hdmi_core_out0_dmareader_rsv_level <= (soc_videooverlaysoc_hdmi_core_out0_dmareader_rsv_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_re) begin
		soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_readable <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_re) begin
			soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_readable <= 1'd0;
		end
	end
	if (((soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_we & soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_writable) & (~soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_replace))) begin
		soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_produce <= (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_produce + 1'd1);
	end
	if (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_do_read) begin
		soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_consume <= (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_we & soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_syncfifo_writable) & (~soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_replace))) begin
		if ((~soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_do_read)) begin
			soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level0 <= (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level0 + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_do_read) begin
			soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level0 <= (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level0 - 1'd1);
		end
	end
	vns_videooutcore_state <= vns_videooutcore_next_state;
	if (soc_videooverlaysoc_hdmi_core_out0_dmareader_offset_next_value_ce) begin
		soc_videooverlaysoc_hdmi_core_out0_dmareader_offset <= soc_videooverlaysoc_hdmi_core_out0_dmareader_offset_next_value;
	end
	soc_videooverlaysoc_hdmi_core_out0_toggle_o_r <= soc_videooverlaysoc_hdmi_core_out0_toggle_o;
	soc_videooverlaysoc_timing_rgb_delay_next_s0 <= soc_videooverlaysoc_timing_rgb_delay_sink_payload_r;
	soc_videooverlaysoc_timing_rgb_delay_next_s1 <= soc_videooverlaysoc_timing_rgb_delay_next_s0;
	soc_videooverlaysoc_timing_rgb_delay_next_s2 <= soc_videooverlaysoc_timing_rgb_delay_next_s1;
	soc_videooverlaysoc_timing_rgb_delay_next_s3 <= soc_videooverlaysoc_timing_rgb_delay_next_s2;
	soc_videooverlaysoc_timing_rgb_delay_next_s4 <= soc_videooverlaysoc_timing_rgb_delay_sink_payload_g;
	soc_videooverlaysoc_timing_rgb_delay_next_s5 <= soc_videooverlaysoc_timing_rgb_delay_next_s4;
	soc_videooverlaysoc_timing_rgb_delay_next_s6 <= soc_videooverlaysoc_timing_rgb_delay_next_s5;
	soc_videooverlaysoc_timing_rgb_delay_next_s7 <= soc_videooverlaysoc_timing_rgb_delay_next_s6;
	soc_videooverlaysoc_timing_rgb_delay_next_s8 <= soc_videooverlaysoc_timing_rgb_delay_sink_payload_b;
	soc_videooverlaysoc_timing_rgb_delay_next_s9 <= soc_videooverlaysoc_timing_rgb_delay_next_s8;
	soc_videooverlaysoc_timing_rgb_delay_next_s10 <= soc_videooverlaysoc_timing_rgb_delay_next_s9;
	soc_videooverlaysoc_timing_rgb_delay_next_s11 <= soc_videooverlaysoc_timing_rgb_delay_next_s10;
	soc_videooverlaysoc_encoder0_n1d <= (((((((soc_videooverlaysoc_encoder0_d0[0] + soc_videooverlaysoc_encoder0_d0[1]) + soc_videooverlaysoc_encoder0_d0[2]) + soc_videooverlaysoc_encoder0_d0[3]) + soc_videooverlaysoc_encoder0_d0[4]) + soc_videooverlaysoc_encoder0_d0[5]) + soc_videooverlaysoc_encoder0_d0[6]) + soc_videooverlaysoc_encoder0_d0[7]);
	soc_videooverlaysoc_encoder0_d1 <= soc_videooverlaysoc_encoder0_d0;
	soc_videooverlaysoc_encoder0_q_m[0] <= soc_videooverlaysoc_encoder0_d1[0];
	soc_videooverlaysoc_encoder0_q_m[1] <= ((soc_videooverlaysoc_encoder0_d1[0] ^ soc_videooverlaysoc_encoder0_d1[1]) ^ soc_videooverlaysoc_encoder0_q_m8_n);
	soc_videooverlaysoc_encoder0_q_m[2] <= ((((soc_videooverlaysoc_encoder0_d1[0] ^ soc_videooverlaysoc_encoder0_d1[1]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[2]) ^ soc_videooverlaysoc_encoder0_q_m8_n);
	soc_videooverlaysoc_encoder0_q_m[3] <= ((((((soc_videooverlaysoc_encoder0_d1[0] ^ soc_videooverlaysoc_encoder0_d1[1]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[2]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[3]) ^ soc_videooverlaysoc_encoder0_q_m8_n);
	soc_videooverlaysoc_encoder0_q_m[4] <= ((((((((soc_videooverlaysoc_encoder0_d1[0] ^ soc_videooverlaysoc_encoder0_d1[1]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[2]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[3]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[4]) ^ soc_videooverlaysoc_encoder0_q_m8_n);
	soc_videooverlaysoc_encoder0_q_m[5] <= ((((((((((soc_videooverlaysoc_encoder0_d1[0] ^ soc_videooverlaysoc_encoder0_d1[1]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[2]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[3]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[4]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[5]) ^ soc_videooverlaysoc_encoder0_q_m8_n);
	soc_videooverlaysoc_encoder0_q_m[6] <= ((((((((((((soc_videooverlaysoc_encoder0_d1[0] ^ soc_videooverlaysoc_encoder0_d1[1]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[2]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[3]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[4]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[5]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[6]) ^ soc_videooverlaysoc_encoder0_q_m8_n);
	soc_videooverlaysoc_encoder0_q_m[7] <= ((((((((((((((soc_videooverlaysoc_encoder0_d1[0] ^ soc_videooverlaysoc_encoder0_d1[1]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[2]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[3]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[4]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[5]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[6]) ^ soc_videooverlaysoc_encoder0_q_m8_n) ^ soc_videooverlaysoc_encoder0_d1[7]) ^ soc_videooverlaysoc_encoder0_q_m8_n);
	soc_videooverlaysoc_encoder0_q_m[8] <= (~soc_videooverlaysoc_encoder0_q_m8_n);
	soc_videooverlaysoc_encoder0_n0q_m <= ((((((((~soc_videooverlaysoc_encoder0_q_m[0]) + (~soc_videooverlaysoc_encoder0_q_m[1])) + (~soc_videooverlaysoc_encoder0_q_m[2])) + (~soc_videooverlaysoc_encoder0_q_m[3])) + (~soc_videooverlaysoc_encoder0_q_m[4])) + (~soc_videooverlaysoc_encoder0_q_m[5])) + (~soc_videooverlaysoc_encoder0_q_m[6])) + (~soc_videooverlaysoc_encoder0_q_m[7]));
	soc_videooverlaysoc_encoder0_n1q_m <= (((((((soc_videooverlaysoc_encoder0_q_m[0] + soc_videooverlaysoc_encoder0_q_m[1]) + soc_videooverlaysoc_encoder0_q_m[2]) + soc_videooverlaysoc_encoder0_q_m[3]) + soc_videooverlaysoc_encoder0_q_m[4]) + soc_videooverlaysoc_encoder0_q_m[5]) + soc_videooverlaysoc_encoder0_q_m[6]) + soc_videooverlaysoc_encoder0_q_m[7]);
	soc_videooverlaysoc_encoder0_q_m_r <= soc_videooverlaysoc_encoder0_q_m;
	soc_videooverlaysoc_encoder0_new_c0 <= soc_videooverlaysoc_encoder0_c;
	soc_videooverlaysoc_encoder0_new_de0 <= soc_videooverlaysoc_encoder0_de;
	soc_videooverlaysoc_encoder0_new_c1 <= soc_videooverlaysoc_encoder0_new_c0;
	soc_videooverlaysoc_encoder0_new_de1 <= soc_videooverlaysoc_encoder0_new_de0;
	soc_videooverlaysoc_encoder0_new_c2 <= soc_videooverlaysoc_encoder0_new_c1;
	soc_videooverlaysoc_encoder0_new_de2 <= soc_videooverlaysoc_encoder0_new_de1;
	if (soc_videooverlaysoc_encoder0_new_de2) begin
		if (((soc_videooverlaysoc_encoder0_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (soc_videooverlaysoc_encoder0_n1q_m == soc_videooverlaysoc_encoder0_n0q_m)}))) begin
			soc_videooverlaysoc_encoder0_out[9] <= (~soc_videooverlaysoc_encoder0_q_m_r[8]);
			soc_videooverlaysoc_encoder0_out[8] <= soc_videooverlaysoc_encoder0_q_m_r[8];
			if (soc_videooverlaysoc_encoder0_q_m_r[8]) begin
				soc_videooverlaysoc_encoder0_out[7:0] <= soc_videooverlaysoc_encoder0_q_m_r[7:0];
				soc_videooverlaysoc_encoder0_cnt <= ((soc_videooverlaysoc_encoder0_cnt + $signed({1'd0, soc_videooverlaysoc_encoder0_n1q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder0_n0q_m}));
			end else begin
				soc_videooverlaysoc_encoder0_out[7:0] <= (~soc_videooverlaysoc_encoder0_q_m_r[7:0]);
				soc_videooverlaysoc_encoder0_cnt <= ((soc_videooverlaysoc_encoder0_cnt + $signed({1'd0, soc_videooverlaysoc_encoder0_n0q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder0_n1q_m}));
			end
		end else begin
			if ((((~soc_videooverlaysoc_encoder0_cnt[5]) & $signed({1'd0, (soc_videooverlaysoc_encoder0_n1q_m > soc_videooverlaysoc_encoder0_n0q_m)})) | (soc_videooverlaysoc_encoder0_cnt[5] & $signed({1'd0, (soc_videooverlaysoc_encoder0_n0q_m > soc_videooverlaysoc_encoder0_n1q_m)})))) begin
				soc_videooverlaysoc_encoder0_out[9] <= 1'd1;
				soc_videooverlaysoc_encoder0_out[8] <= soc_videooverlaysoc_encoder0_q_m_r[8];
				soc_videooverlaysoc_encoder0_out[7:0] <= (~soc_videooverlaysoc_encoder0_q_m_r[7:0]);
				soc_videooverlaysoc_encoder0_cnt <= (((soc_videooverlaysoc_encoder0_cnt + $signed({1'd0, {soc_videooverlaysoc_encoder0_q_m_r[8], 1'd0}})) + $signed({1'd0, soc_videooverlaysoc_encoder0_n0q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder0_n1q_m}));
			end else begin
				soc_videooverlaysoc_encoder0_out[9] <= 1'd0;
				soc_videooverlaysoc_encoder0_out[8] <= soc_videooverlaysoc_encoder0_q_m_r[8];
				soc_videooverlaysoc_encoder0_out[7:0] <= soc_videooverlaysoc_encoder0_q_m_r[7:0];
				soc_videooverlaysoc_encoder0_cnt <= (((soc_videooverlaysoc_encoder0_cnt - $signed({1'd0, {(~soc_videooverlaysoc_encoder0_q_m_r[8]), 1'd0}})) + $signed({1'd0, soc_videooverlaysoc_encoder0_n1q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder0_n0q_m}));
			end
		end
	end else begin
		soc_videooverlaysoc_encoder0_out <= vns_sync_f_array_muxed0;
		soc_videooverlaysoc_encoder0_cnt <= 1'd0;
	end
	soc_videooverlaysoc_encoder1_n1d <= (((((((soc_videooverlaysoc_encoder1_d0[0] + soc_videooverlaysoc_encoder1_d0[1]) + soc_videooverlaysoc_encoder1_d0[2]) + soc_videooverlaysoc_encoder1_d0[3]) + soc_videooverlaysoc_encoder1_d0[4]) + soc_videooverlaysoc_encoder1_d0[5]) + soc_videooverlaysoc_encoder1_d0[6]) + soc_videooverlaysoc_encoder1_d0[7]);
	soc_videooverlaysoc_encoder1_d1 <= soc_videooverlaysoc_encoder1_d0;
	soc_videooverlaysoc_encoder1_q_m[0] <= soc_videooverlaysoc_encoder1_d1[0];
	soc_videooverlaysoc_encoder1_q_m[1] <= ((soc_videooverlaysoc_encoder1_d1[0] ^ soc_videooverlaysoc_encoder1_d1[1]) ^ soc_videooverlaysoc_encoder1_q_m8_n);
	soc_videooverlaysoc_encoder1_q_m[2] <= ((((soc_videooverlaysoc_encoder1_d1[0] ^ soc_videooverlaysoc_encoder1_d1[1]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[2]) ^ soc_videooverlaysoc_encoder1_q_m8_n);
	soc_videooverlaysoc_encoder1_q_m[3] <= ((((((soc_videooverlaysoc_encoder1_d1[0] ^ soc_videooverlaysoc_encoder1_d1[1]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[2]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[3]) ^ soc_videooverlaysoc_encoder1_q_m8_n);
	soc_videooverlaysoc_encoder1_q_m[4] <= ((((((((soc_videooverlaysoc_encoder1_d1[0] ^ soc_videooverlaysoc_encoder1_d1[1]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[2]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[3]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[4]) ^ soc_videooverlaysoc_encoder1_q_m8_n);
	soc_videooverlaysoc_encoder1_q_m[5] <= ((((((((((soc_videooverlaysoc_encoder1_d1[0] ^ soc_videooverlaysoc_encoder1_d1[1]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[2]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[3]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[4]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[5]) ^ soc_videooverlaysoc_encoder1_q_m8_n);
	soc_videooverlaysoc_encoder1_q_m[6] <= ((((((((((((soc_videooverlaysoc_encoder1_d1[0] ^ soc_videooverlaysoc_encoder1_d1[1]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[2]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[3]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[4]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[5]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[6]) ^ soc_videooverlaysoc_encoder1_q_m8_n);
	soc_videooverlaysoc_encoder1_q_m[7] <= ((((((((((((((soc_videooverlaysoc_encoder1_d1[0] ^ soc_videooverlaysoc_encoder1_d1[1]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[2]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[3]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[4]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[5]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[6]) ^ soc_videooverlaysoc_encoder1_q_m8_n) ^ soc_videooverlaysoc_encoder1_d1[7]) ^ soc_videooverlaysoc_encoder1_q_m8_n);
	soc_videooverlaysoc_encoder1_q_m[8] <= (~soc_videooverlaysoc_encoder1_q_m8_n);
	soc_videooverlaysoc_encoder1_n0q_m <= ((((((((~soc_videooverlaysoc_encoder1_q_m[0]) + (~soc_videooverlaysoc_encoder1_q_m[1])) + (~soc_videooverlaysoc_encoder1_q_m[2])) + (~soc_videooverlaysoc_encoder1_q_m[3])) + (~soc_videooverlaysoc_encoder1_q_m[4])) + (~soc_videooverlaysoc_encoder1_q_m[5])) + (~soc_videooverlaysoc_encoder1_q_m[6])) + (~soc_videooverlaysoc_encoder1_q_m[7]));
	soc_videooverlaysoc_encoder1_n1q_m <= (((((((soc_videooverlaysoc_encoder1_q_m[0] + soc_videooverlaysoc_encoder1_q_m[1]) + soc_videooverlaysoc_encoder1_q_m[2]) + soc_videooverlaysoc_encoder1_q_m[3]) + soc_videooverlaysoc_encoder1_q_m[4]) + soc_videooverlaysoc_encoder1_q_m[5]) + soc_videooverlaysoc_encoder1_q_m[6]) + soc_videooverlaysoc_encoder1_q_m[7]);
	soc_videooverlaysoc_encoder1_q_m_r <= soc_videooverlaysoc_encoder1_q_m;
	soc_videooverlaysoc_encoder1_new_c0 <= soc_videooverlaysoc_encoder1_c;
	soc_videooverlaysoc_encoder1_new_de0 <= soc_videooverlaysoc_encoder1_de;
	soc_videooverlaysoc_encoder1_new_c1 <= soc_videooverlaysoc_encoder1_new_c0;
	soc_videooverlaysoc_encoder1_new_de1 <= soc_videooverlaysoc_encoder1_new_de0;
	soc_videooverlaysoc_encoder1_new_c2 <= soc_videooverlaysoc_encoder1_new_c1;
	soc_videooverlaysoc_encoder1_new_de2 <= soc_videooverlaysoc_encoder1_new_de1;
	if (soc_videooverlaysoc_encoder1_new_de2) begin
		if (((soc_videooverlaysoc_encoder1_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (soc_videooverlaysoc_encoder1_n1q_m == soc_videooverlaysoc_encoder1_n0q_m)}))) begin
			soc_videooverlaysoc_encoder1_out[9] <= (~soc_videooverlaysoc_encoder1_q_m_r[8]);
			soc_videooverlaysoc_encoder1_out[8] <= soc_videooverlaysoc_encoder1_q_m_r[8];
			if (soc_videooverlaysoc_encoder1_q_m_r[8]) begin
				soc_videooverlaysoc_encoder1_out[7:0] <= soc_videooverlaysoc_encoder1_q_m_r[7:0];
				soc_videooverlaysoc_encoder1_cnt <= ((soc_videooverlaysoc_encoder1_cnt + $signed({1'd0, soc_videooverlaysoc_encoder1_n1q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder1_n0q_m}));
			end else begin
				soc_videooverlaysoc_encoder1_out[7:0] <= (~soc_videooverlaysoc_encoder1_q_m_r[7:0]);
				soc_videooverlaysoc_encoder1_cnt <= ((soc_videooverlaysoc_encoder1_cnt + $signed({1'd0, soc_videooverlaysoc_encoder1_n0q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder1_n1q_m}));
			end
		end else begin
			if ((((~soc_videooverlaysoc_encoder1_cnt[5]) & $signed({1'd0, (soc_videooverlaysoc_encoder1_n1q_m > soc_videooverlaysoc_encoder1_n0q_m)})) | (soc_videooverlaysoc_encoder1_cnt[5] & $signed({1'd0, (soc_videooverlaysoc_encoder1_n0q_m > soc_videooverlaysoc_encoder1_n1q_m)})))) begin
				soc_videooverlaysoc_encoder1_out[9] <= 1'd1;
				soc_videooverlaysoc_encoder1_out[8] <= soc_videooverlaysoc_encoder1_q_m_r[8];
				soc_videooverlaysoc_encoder1_out[7:0] <= (~soc_videooverlaysoc_encoder1_q_m_r[7:0]);
				soc_videooverlaysoc_encoder1_cnt <= (((soc_videooverlaysoc_encoder1_cnt + $signed({1'd0, {soc_videooverlaysoc_encoder1_q_m_r[8], 1'd0}})) + $signed({1'd0, soc_videooverlaysoc_encoder1_n0q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder1_n1q_m}));
			end else begin
				soc_videooverlaysoc_encoder1_out[9] <= 1'd0;
				soc_videooverlaysoc_encoder1_out[8] <= soc_videooverlaysoc_encoder1_q_m_r[8];
				soc_videooverlaysoc_encoder1_out[7:0] <= soc_videooverlaysoc_encoder1_q_m_r[7:0];
				soc_videooverlaysoc_encoder1_cnt <= (((soc_videooverlaysoc_encoder1_cnt - $signed({1'd0, {(~soc_videooverlaysoc_encoder1_q_m_r[8]), 1'd0}})) + $signed({1'd0, soc_videooverlaysoc_encoder1_n1q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder1_n0q_m}));
			end
		end
	end else begin
		soc_videooverlaysoc_encoder1_out <= vns_sync_f_array_muxed1;
		soc_videooverlaysoc_encoder1_cnt <= 1'd0;
	end
	soc_videooverlaysoc_encoder2_n1d <= (((((((soc_videooverlaysoc_encoder2_d0[0] + soc_videooverlaysoc_encoder2_d0[1]) + soc_videooverlaysoc_encoder2_d0[2]) + soc_videooverlaysoc_encoder2_d0[3]) + soc_videooverlaysoc_encoder2_d0[4]) + soc_videooverlaysoc_encoder2_d0[5]) + soc_videooverlaysoc_encoder2_d0[6]) + soc_videooverlaysoc_encoder2_d0[7]);
	soc_videooverlaysoc_encoder2_d1 <= soc_videooverlaysoc_encoder2_d0;
	soc_videooverlaysoc_encoder2_q_m[0] <= soc_videooverlaysoc_encoder2_d1[0];
	soc_videooverlaysoc_encoder2_q_m[1] <= ((soc_videooverlaysoc_encoder2_d1[0] ^ soc_videooverlaysoc_encoder2_d1[1]) ^ soc_videooverlaysoc_encoder2_q_m8_n);
	soc_videooverlaysoc_encoder2_q_m[2] <= ((((soc_videooverlaysoc_encoder2_d1[0] ^ soc_videooverlaysoc_encoder2_d1[1]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[2]) ^ soc_videooverlaysoc_encoder2_q_m8_n);
	soc_videooverlaysoc_encoder2_q_m[3] <= ((((((soc_videooverlaysoc_encoder2_d1[0] ^ soc_videooverlaysoc_encoder2_d1[1]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[2]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[3]) ^ soc_videooverlaysoc_encoder2_q_m8_n);
	soc_videooverlaysoc_encoder2_q_m[4] <= ((((((((soc_videooverlaysoc_encoder2_d1[0] ^ soc_videooverlaysoc_encoder2_d1[1]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[2]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[3]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[4]) ^ soc_videooverlaysoc_encoder2_q_m8_n);
	soc_videooverlaysoc_encoder2_q_m[5] <= ((((((((((soc_videooverlaysoc_encoder2_d1[0] ^ soc_videooverlaysoc_encoder2_d1[1]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[2]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[3]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[4]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[5]) ^ soc_videooverlaysoc_encoder2_q_m8_n);
	soc_videooverlaysoc_encoder2_q_m[6] <= ((((((((((((soc_videooverlaysoc_encoder2_d1[0] ^ soc_videooverlaysoc_encoder2_d1[1]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[2]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[3]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[4]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[5]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[6]) ^ soc_videooverlaysoc_encoder2_q_m8_n);
	soc_videooverlaysoc_encoder2_q_m[7] <= ((((((((((((((soc_videooverlaysoc_encoder2_d1[0] ^ soc_videooverlaysoc_encoder2_d1[1]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[2]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[3]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[4]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[5]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[6]) ^ soc_videooverlaysoc_encoder2_q_m8_n) ^ soc_videooverlaysoc_encoder2_d1[7]) ^ soc_videooverlaysoc_encoder2_q_m8_n);
	soc_videooverlaysoc_encoder2_q_m[8] <= (~soc_videooverlaysoc_encoder2_q_m8_n);
	soc_videooverlaysoc_encoder2_n0q_m <= ((((((((~soc_videooverlaysoc_encoder2_q_m[0]) + (~soc_videooverlaysoc_encoder2_q_m[1])) + (~soc_videooverlaysoc_encoder2_q_m[2])) + (~soc_videooverlaysoc_encoder2_q_m[3])) + (~soc_videooverlaysoc_encoder2_q_m[4])) + (~soc_videooverlaysoc_encoder2_q_m[5])) + (~soc_videooverlaysoc_encoder2_q_m[6])) + (~soc_videooverlaysoc_encoder2_q_m[7]));
	soc_videooverlaysoc_encoder2_n1q_m <= (((((((soc_videooverlaysoc_encoder2_q_m[0] + soc_videooverlaysoc_encoder2_q_m[1]) + soc_videooverlaysoc_encoder2_q_m[2]) + soc_videooverlaysoc_encoder2_q_m[3]) + soc_videooverlaysoc_encoder2_q_m[4]) + soc_videooverlaysoc_encoder2_q_m[5]) + soc_videooverlaysoc_encoder2_q_m[6]) + soc_videooverlaysoc_encoder2_q_m[7]);
	soc_videooverlaysoc_encoder2_q_m_r <= soc_videooverlaysoc_encoder2_q_m;
	soc_videooverlaysoc_encoder2_new_c0 <= soc_videooverlaysoc_encoder2_c;
	soc_videooverlaysoc_encoder2_new_de0 <= soc_videooverlaysoc_encoder2_de;
	soc_videooverlaysoc_encoder2_new_c1 <= soc_videooverlaysoc_encoder2_new_c0;
	soc_videooverlaysoc_encoder2_new_de1 <= soc_videooverlaysoc_encoder2_new_de0;
	soc_videooverlaysoc_encoder2_new_c2 <= soc_videooverlaysoc_encoder2_new_c1;
	soc_videooverlaysoc_encoder2_new_de2 <= soc_videooverlaysoc_encoder2_new_de1;
	if (soc_videooverlaysoc_encoder2_new_de2) begin
		if (((soc_videooverlaysoc_encoder2_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (soc_videooverlaysoc_encoder2_n1q_m == soc_videooverlaysoc_encoder2_n0q_m)}))) begin
			soc_videooverlaysoc_encoder2_out[9] <= (~soc_videooverlaysoc_encoder2_q_m_r[8]);
			soc_videooverlaysoc_encoder2_out[8] <= soc_videooverlaysoc_encoder2_q_m_r[8];
			if (soc_videooverlaysoc_encoder2_q_m_r[8]) begin
				soc_videooverlaysoc_encoder2_out[7:0] <= soc_videooverlaysoc_encoder2_q_m_r[7:0];
				soc_videooverlaysoc_encoder2_cnt <= ((soc_videooverlaysoc_encoder2_cnt + $signed({1'd0, soc_videooverlaysoc_encoder2_n1q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder2_n0q_m}));
			end else begin
				soc_videooverlaysoc_encoder2_out[7:0] <= (~soc_videooverlaysoc_encoder2_q_m_r[7:0]);
				soc_videooverlaysoc_encoder2_cnt <= ((soc_videooverlaysoc_encoder2_cnt + $signed({1'd0, soc_videooverlaysoc_encoder2_n0q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder2_n1q_m}));
			end
		end else begin
			if ((((~soc_videooverlaysoc_encoder2_cnt[5]) & $signed({1'd0, (soc_videooverlaysoc_encoder2_n1q_m > soc_videooverlaysoc_encoder2_n0q_m)})) | (soc_videooverlaysoc_encoder2_cnt[5] & $signed({1'd0, (soc_videooverlaysoc_encoder2_n0q_m > soc_videooverlaysoc_encoder2_n1q_m)})))) begin
				soc_videooverlaysoc_encoder2_out[9] <= 1'd1;
				soc_videooverlaysoc_encoder2_out[8] <= soc_videooverlaysoc_encoder2_q_m_r[8];
				soc_videooverlaysoc_encoder2_out[7:0] <= (~soc_videooverlaysoc_encoder2_q_m_r[7:0]);
				soc_videooverlaysoc_encoder2_cnt <= (((soc_videooverlaysoc_encoder2_cnt + $signed({1'd0, {soc_videooverlaysoc_encoder2_q_m_r[8], 1'd0}})) + $signed({1'd0, soc_videooverlaysoc_encoder2_n0q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder2_n1q_m}));
			end else begin
				soc_videooverlaysoc_encoder2_out[9] <= 1'd0;
				soc_videooverlaysoc_encoder2_out[8] <= soc_videooverlaysoc_encoder2_q_m_r[8];
				soc_videooverlaysoc_encoder2_out[7:0] <= soc_videooverlaysoc_encoder2_q_m_r[7:0];
				soc_videooverlaysoc_encoder2_cnt <= (((soc_videooverlaysoc_encoder2_cnt - $signed({1'd0, {(~soc_videooverlaysoc_encoder2_q_m_r[8]), 1'd0}})) + $signed({1'd0, soc_videooverlaysoc_encoder2_n1q_m})) - $signed({1'd0, soc_videooverlaysoc_encoder2_n0q_m}));
			end
		end
	end else begin
		soc_videooverlaysoc_encoder2_out <= vns_sync_f_array_muxed2;
		soc_videooverlaysoc_encoder2_cnt <= 1'd0;
	end
	soc_videooverlaysoc_in0_de <= soc_videooverlaysoc_hdmi_in0_timing_payload_de;
	soc_videooverlaysoc_in0_de_r <= soc_videooverlaysoc_in0_de;
	soc_videooverlaysoc_in0_vsync <= soc_videooverlaysoc_hdmi_in0_timing_payload_vsync;
	soc_videooverlaysoc_in0_vsync_r <= soc_videooverlaysoc_in0_vsync;
	soc_videooverlaysoc_in0_hsync <= soc_videooverlaysoc_hdmi_in0_timing_payload_hsync;
	soc_videooverlaysoc_in0_hsync_r <= soc_videooverlaysoc_in0_hsync;
	if ((soc_videooverlaysoc_in0_vsync & (~soc_videooverlaysoc_in0_vsync_r))) begin
		soc_videooverlaysoc_vcounter <= 1'd0;
	end else begin
		if ((soc_videooverlaysoc_in0_de & (~soc_videooverlaysoc_in0_de_r))) begin
			soc_videooverlaysoc_vcounter <= (soc_videooverlaysoc_vcounter + 1'd1);
		end
	end
	if ((soc_videooverlaysoc_in0_de & (~soc_videooverlaysoc_in0_de_r))) begin
		soc_videooverlaysoc_hcounter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_in0_de) begin
			soc_videooverlaysoc_hcounter <= (soc_videooverlaysoc_hcounter + 1'd1);
		end
	end
	if (pix_o_rst) begin
		soc_videooverlaysoc_hdmi_in0_syncpol_c0 <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_syncpol_c1 <= 10'd0;
		soc_videooverlaysoc_hdmi_in0_syncpol_c2 <= 10'd0;
		soc_videooverlaysoc_hdmi_out0_clk_gen_ce <= 1'd0;
		soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c0 <= 10'd0;
		soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c1 <= 10'd0;
		soc_videooverlaysoc_hdmi_out0_phy_sink_payload_c2 <= 11'd0;
		soc_videooverlaysoc_hdmi_out0_phy_es0_ce <= 1'd0;
		soc_videooverlaysoc_hdmi_out0_phy_es1_ce <= 1'd0;
		soc_videooverlaysoc_hdmi_out0_phy_es2_ce <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_timing_valid <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_timing_payload_hsync <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_timing_payload_vsync <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_timing_payload_de <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_syncpol_c0 <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_syncpol_c1 <= 10'd0;
		soc_videooverlaysoc_hdmi_in1_syncpol_c2 <= 10'd0;
		soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q <= 3'd0;
		soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q_binary <= 3'd0;
		soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q <= 5'd0;
		soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q_binary <= 5'd0;
		soc_videooverlaysoc_out_dram_port_cmd_buffer_level <= 3'd0;
		soc_videooverlaysoc_out_dram_port_cmd_buffer_produce <= 2'd0;
		soc_videooverlaysoc_out_dram_port_cmd_buffer_consume <= 2'd0;
		soc_videooverlaysoc_out_dram_port_counter <= 3'd0;
		soc_videooverlaysoc_out_dram_port_rdata_buffer_source_payload_data <= 256'd0;
		soc_videooverlaysoc_out_dram_port_rdata_buffer_valid_n <= 1'd0;
		soc_videooverlaysoc_out_dram_port_rdata_buffer_first_n <= 1'd0;
		soc_videooverlaysoc_out_dram_port_rdata_buffer_last_n <= 1'd0;
		soc_videooverlaysoc_out_dram_port_rdata_converter_converter_mux <= 3'd0;
		soc_videooverlaysoc_out_dram_port_rdata_chunk <= 8'd1;
		soc_videooverlaysoc_hdmi_core_out0_underflow_counter_status <= 32'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q <= 2'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q_binary <= 2'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_rsv_level <= 11'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_readable <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_level0 <= 11'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_produce <= 10'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_consume <= 10'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_offset <= 27'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_v <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_v_r <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_sof <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_underflow_counter <= 32'd0;
		soc_videooverlaysoc_core_source_valid_d <= 1'd0;
		soc_videooverlaysoc_core_source_data_d <= 32'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s0 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s1 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s2 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s3 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s4 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s5 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s6 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s7 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s8 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s9 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s10 <= 8'd0;
		soc_videooverlaysoc_timing_rgb_delay_next_s11 <= 8'd0;
		soc_videooverlaysoc_hdcp_hpd <= 1'd0;
		soc_videooverlaysoc_hdcp_hdcp_ena <= 1'd0;
		soc_videooverlaysoc_hdcp_Aksv14_write <= 1'd0;
		soc_videooverlaysoc_hdcp_ctl_code <= 4'd0;
		soc_videooverlaysoc_hdcp_An <= 64'd0;
		soc_videooverlaysoc_Aksv14_r <= 1'd0;
		soc_videooverlaysoc_encoder0_out <= 10'd0;
		soc_videooverlaysoc_encoder0_d1 <= 8'd0;
		soc_videooverlaysoc_encoder0_n1d <= 4'd0;
		soc_videooverlaysoc_encoder0_q_m <= 9'd0;
		soc_videooverlaysoc_encoder0_q_m_r <= 9'd0;
		soc_videooverlaysoc_encoder0_n0q_m <= 4'd0;
		soc_videooverlaysoc_encoder0_n1q_m <= 4'd0;
		soc_videooverlaysoc_encoder0_cnt <= 6'sd64;
		soc_videooverlaysoc_encoder0_new_c0 <= 2'd0;
		soc_videooverlaysoc_encoder0_new_de0 <= 1'd0;
		soc_videooverlaysoc_encoder0_new_c1 <= 2'd0;
		soc_videooverlaysoc_encoder0_new_de1 <= 1'd0;
		soc_videooverlaysoc_encoder0_new_c2 <= 2'd0;
		soc_videooverlaysoc_encoder0_new_de2 <= 1'd0;
		soc_videooverlaysoc_encoder1_out <= 10'd0;
		soc_videooverlaysoc_encoder1_d1 <= 8'd0;
		soc_videooverlaysoc_encoder1_n1d <= 4'd0;
		soc_videooverlaysoc_encoder1_q_m <= 9'd0;
		soc_videooverlaysoc_encoder1_q_m_r <= 9'd0;
		soc_videooverlaysoc_encoder1_n0q_m <= 4'd0;
		soc_videooverlaysoc_encoder1_n1q_m <= 4'd0;
		soc_videooverlaysoc_encoder1_cnt <= 6'sd64;
		soc_videooverlaysoc_encoder1_new_c0 <= 2'd0;
		soc_videooverlaysoc_encoder1_new_de0 <= 1'd0;
		soc_videooverlaysoc_encoder1_new_c1 <= 2'd0;
		soc_videooverlaysoc_encoder1_new_de1 <= 1'd0;
		soc_videooverlaysoc_encoder1_new_c2 <= 2'd0;
		soc_videooverlaysoc_encoder1_new_de2 <= 1'd0;
		soc_videooverlaysoc_encoder2_out <= 10'd0;
		soc_videooverlaysoc_encoder2_d1 <= 8'd0;
		soc_videooverlaysoc_encoder2_n1d <= 4'd0;
		soc_videooverlaysoc_encoder2_q_m <= 9'd0;
		soc_videooverlaysoc_encoder2_q_m_r <= 9'd0;
		soc_videooverlaysoc_encoder2_n0q_m <= 4'd0;
		soc_videooverlaysoc_encoder2_n1q_m <= 4'd0;
		soc_videooverlaysoc_encoder2_cnt <= 6'sd64;
		soc_videooverlaysoc_encoder2_new_c0 <= 2'd0;
		soc_videooverlaysoc_encoder2_new_de0 <= 1'd0;
		soc_videooverlaysoc_encoder2_new_c1 <= 2'd0;
		soc_videooverlaysoc_encoder2_new_de1 <= 1'd0;
		soc_videooverlaysoc_encoder2_new_c2 <= 2'd0;
		soc_videooverlaysoc_encoder2_new_de2 <= 1'd0;
		soc_videooverlaysoc_c0_pix_o <= 10'd0;
		soc_videooverlaysoc_c1_pix_o <= 10'd0;
		soc_videooverlaysoc_c2_pix_o <= 10'd0;
		soc_videooverlaysoc_c0_next0 <= 10'd0;
		soc_videooverlaysoc_c1_next0 <= 10'd0;
		soc_videooverlaysoc_c2_next0 <= 10'd0;
		soc_videooverlaysoc_c0_next1 <= 10'd0;
		soc_videooverlaysoc_c1_next1 <= 10'd0;
		soc_videooverlaysoc_c2_next1 <= 10'd0;
		soc_videooverlaysoc_c0_next2 <= 10'd0;
		soc_videooverlaysoc_c1_next2 <= 10'd0;
		soc_videooverlaysoc_c2_next2 <= 10'd0;
		soc_videooverlaysoc_c0_next3 <= 10'd0;
		soc_videooverlaysoc_c1_next3 <= 10'd0;
		soc_videooverlaysoc_c2_next3 <= 10'd0;
		soc_videooverlaysoc_c0_next4 <= 10'd0;
		soc_videooverlaysoc_c1_next4 <= 10'd0;
		soc_videooverlaysoc_c2_next4 <= 10'd0;
		soc_videooverlaysoc_c0_next5 <= 10'd0;
		soc_videooverlaysoc_c1_next5 <= 10'd0;
		soc_videooverlaysoc_c2_next5 <= 10'd0;
		soc_videooverlaysoc_hcounter <= 12'd0;
		soc_videooverlaysoc_vcounter <= 12'd0;
		soc_videooverlaysoc_in0_de <= 1'd0;
		soc_videooverlaysoc_in0_de_r <= 1'd0;
		soc_videooverlaysoc_in0_vsync <= 1'd0;
		soc_videooverlaysoc_in0_vsync_r <= 1'd0;
		soc_videooverlaysoc_in0_hsync <= 1'd0;
		soc_videooverlaysoc_in0_hsync_r <= 1'd0;
		vns_videooutcore_state <= 2'd0;
	end
	vns_xilinxmultiregimpl84_regs0 <= soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q;
	vns_xilinxmultiregimpl84_regs1 <= vns_xilinxmultiregimpl84_regs0;
	vns_xilinxmultiregimpl85_regs0 <= soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q;
	vns_xilinxmultiregimpl85_regs1 <= vns_xilinxmultiregimpl85_regs0;
	vns_xilinxmultiregimpl87_regs0 <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q;
	vns_xilinxmultiregimpl87_regs1 <= vns_xilinxmultiregimpl87_regs0;
	vns_xilinxmultiregimpl90_regs0 <= soc_videooverlaysoc_hdmi_core_out0_toggle_i;
	vns_xilinxmultiregimpl90_regs1 <= vns_xilinxmultiregimpl90_regs0;
	vns_xilinxmultiregimpl91_regs0 <= soc_videooverlaysoc_i2c_snoop_Aksv14_write;
	vns_xilinxmultiregimpl91_regs1 <= vns_xilinxmultiregimpl91_regs0;
end

always @(posedge sys_clk) begin
	soc_videooverlaysoc_videooverlaysoc_sys_counter <= (soc_videooverlaysoc_videooverlaysoc_sys_counter + 1'd1);
	fpga_led40 <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors != 32'd4294967295)) begin
		if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_error) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors + 1'd1);
		end
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_o_rsp_data;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_cpu_reset <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_reset_debug_logic | sys_rst);
	if (((((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_stb & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_cyc) & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_in_progress)) & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_complete)) & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_wait_for_ack))) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_data <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_dat_w;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_address <= ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_adr[5:0] <<< 2'd2) | 1'd0);
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_wr <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_we;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_valid <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_in_progress <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_complete <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_ack <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_in_progress) begin
			if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_o_cmd_ready) begin
				soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_valid <= 1'd0;
				soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_wr <= 1'd0;
				soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_complete <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_in_progress <= 1'd0;
			end
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_complete) begin
				soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_complete <= 1'd0;
				soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_ack <= 1'd1;
				soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_wait_for_ack <= 1'd1;
			end else begin
				if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_wait_for_ack & (~(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_stb & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_cyc)))) begin
					soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_wait_for_ack <= 1'd0;
					soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_ack <= 1'd0;
				end
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_o_resetOut) begin
		if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_cyc & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_stb)) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_err <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_err <= 1'd0;
		end
		if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_cyc & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_stb)) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_d_err <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_d_err <= 1'd0;
		end
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_reset_debug_logic <= 1'd1;
	end else begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_reset_debug_logic <= 1'd0;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_ack <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_cyc & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_stb) & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_ack))) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_ack <= 1'd1;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_ack <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_cyc & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_stb) & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_ack))) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_ack <= 1'd1;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_dat_w;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_adr;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_dat_r <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_r;
	if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_counter == 1'd1)) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_we;
	end
	if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_counter == 2'd2)) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_ack <= 1'd1;
	end
	if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_counter == 2'd3)) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_ack <= 1'd0;
	end
	if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_counter != 1'd0)) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_counter <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_counter + 1'd1);
	end else begin
		if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_cyc & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_stb)) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_counter <= 1'd1;
		end
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_ready <= 1'd0;
	if (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_valid & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_busy)) & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_ready))) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_reg <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_payload_data;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_bitcount <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_busy <= 1'd1;
		serial_tx <= 1'd0;
	end else begin
		if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_uart_clk_txen & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_busy)) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_bitcount <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_bitcount + 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_bitcount == 4'd8)) begin
				serial_tx <= 1'd1;
			end else begin
				if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_bitcount == 4'd9)) begin
					serial_tx <= 1'd1;
					soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_busy <= 1'd0;
					soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_ready <= 1'd1;
				end else begin
					serial_tx <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_reg[0];
					soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_reg <= {1'd0, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_reg[7:1]};
				end
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_busy) begin
		{soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_uart_clk_txen, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_phase_accumulator_tx} <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_phase_accumulator_tx + soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage);
	end else begin
		{soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_uart_clk_txen, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_phase_accumulator_tx} <= 1'd0;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_valid <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_r <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx;
	if ((~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_busy)) begin
		if (((~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_r)) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_busy <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_bitcount <= 1'd0;
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_uart_clk_rxen) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_bitcount <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_bitcount + 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_bitcount == 1'd0)) begin
				if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx) begin
					soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_busy <= 1'd0;
				end
			end else begin
				if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_bitcount == 4'd9)) begin
					soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_busy <= 1'd0;
					if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx) begin
						soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_payload_data <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_reg;
						soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_valid <= 1'd1;
					end
				end else begin
					soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_reg <= {soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_reg[7:1]};
				end
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_busy) begin
		{soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_uart_clk_rxen, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_phase_accumulator_rx} <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_phase_accumulator_rx + soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage);
	end else begin
		{soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_uart_clk_rxen, soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_phase_accumulator_rx} <= 32'd2147483648;
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_clear) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_pending <= 1'd0;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_old_trigger <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_trigger;
	if (((~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_trigger) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_old_trigger)) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_pending <= 1'd1;
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_clear) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_pending <= 1'd0;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_old_trigger <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_trigger;
	if (((~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_trigger) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_old_trigger)) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_pending <= 1'd1;
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_readable <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_re) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_readable <= 1'd0;
		end
	end
	if (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_we & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_writable) & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_replace))) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_produce <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_produce + 1'd1);
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_do_read) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_consume <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_we & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_syncfifo_writable) & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_replace))) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_do_read)) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level0 <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level0 + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_do_read) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level0 <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level0 - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_readable <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_re) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_readable <= 1'd0;
		end
	end
	if (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_we & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_writable) & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_replace))) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_produce <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_produce + 1'd1);
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_do_read) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_consume <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_we & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_syncfifo_writable) & (~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_replace))) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_do_read)) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level0 <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level0 + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_do_read) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level0 <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level0 - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_reset) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_pending <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_old_trigger <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_pending <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_old_trigger <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_readable <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level0 <= 5'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_produce <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_consume <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_readable <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level0 <= 5'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_produce <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_consume <= 4'd0;
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_storage) begin
		if ((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value == 1'd0)) begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value <= (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value - 1'd1);
		end
	end else begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage;
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_update_value_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value_status <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value;
	end
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_clear) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_pending <= 1'd0;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_old_trigger <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_trigger;
	if (((~soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_trigger) & soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_old_trigger)) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_pending <= 1'd1;
	end
	if (soc_videooverlaysoc_videooverlaysoc_drdy) begin
		case (soc_videooverlaysoc_videooverlaysoc_channel)
			1'd0: begin
				soc_videooverlaysoc_videooverlaysoc_temperature_status <= (soc_videooverlaysoc_videooverlaysoc_data >>> 3'd4);
			end
			1'd1: begin
				soc_videooverlaysoc_videooverlaysoc_vccint_status <= (soc_videooverlaysoc_videooverlaysoc_data >>> 3'd4);
			end
			2'd2: begin
				soc_videooverlaysoc_videooverlaysoc_vccaux_status <= (soc_videooverlaysoc_videooverlaysoc_data >>> 3'd4);
			end
			3'd6: begin
				soc_videooverlaysoc_videooverlaysoc_vccbram_status <= (soc_videooverlaysoc_videooverlaysoc_data >>> 3'd4);
			end
		endcase
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_value + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3]) begin
		if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_value <= 1'd0;
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_re) begin
				soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_value <= (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_value + 1'd1);
			end
		end
	end
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en0 <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata_en;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en1 <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en0;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en2 <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en1;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en3 <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en2;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en4 <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en3;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en5 <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en4;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en6 <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en5;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en7 <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en6;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en7;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en7;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en7;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata_valid <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en7;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en[2:0], soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_en};
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dqs <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe;
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r[14:7];
		end
	endcase
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r <= {soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_i, soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r[15:8]};
	case (soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_value)
		1'd0: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r[7:0];
		end
		1'd1: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r[8:1];
		end
		2'd2: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r[9:2];
		end
		2'd3: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r[10:3];
		end
		3'd4: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r[11:4];
		end
		3'd5: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r[12:5];
		end
		3'd6: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r[13:6];
		end
		3'd7: begin
			soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r[14:7];
		end
	endcase
	if (soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p0_rddata;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p1_rddata;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p2_rddata;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status <= soc_videooverlaysoc_videooverlaysoc_sdram_inti_p3_rddata;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_a <= 11'd1024;
	soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ba <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_cas <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ras <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_we <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_seq_done <= 1'd0;
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_counter == 1'd1)) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ras <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_we <= 1'd1;
	end
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_counter == 3'd4)) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_cas <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ras <= 1'd1;
	end
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_counter == 5'd18)) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_seq_done <= 1'd1;
	end
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_counter == 5'd18)) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_counter <= 1'd0;
	end else begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_counter != 1'd0)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_counter <= (soc_videooverlaysoc_videooverlaysoc_sdram_counter + 1'd1);
		end else begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_seq_start) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_counter <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_wait) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_done)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_count - 1'd1);
		end
	end else begin
		soc_videooverlaysoc_videooverlaysoc_sdram_count <= 10'd782;
	end
	vns_refresher_state <= vns_refresher_next_state;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_close) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_opened <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_open) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_opened <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_replace))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_produce <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_do_read) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_consume <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_replace))) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_do_read)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_do_read) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_valid_n <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_valid;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_first_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_first);
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_last_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_last);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_we <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_payload_we;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_addr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_sink_payload_addr;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_count <= 3'd4;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_ready <= 1'd1;
			end
		end
	end
	vns_bankmachine0_state <= vns_bankmachine0_next_state;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_close) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_opened <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_open) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_opened <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_replace))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_produce <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_do_read) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_consume <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_replace))) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_do_read)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_do_read) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_valid_n <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_valid;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_first_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_first);
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_last_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_last);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_we <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_payload_we;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_addr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_sink_payload_addr;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_count <= 3'd4;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_ready <= 1'd1;
			end
		end
	end
	vns_bankmachine1_state <= vns_bankmachine1_next_state;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_close) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_opened <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_open) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_opened <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_replace))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_produce <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_do_read) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_consume <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_replace))) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_do_read)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_do_read) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_valid_n <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_valid;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_first_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_first);
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_last_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_last);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_we <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_payload_we;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_addr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_sink_payload_addr;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_count <= 3'd4;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_ready <= 1'd1;
			end
		end
	end
	vns_bankmachine2_state <= vns_bankmachine2_next_state;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_close) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_opened <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_open) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_opened <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_replace))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_produce <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_do_read) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_consume <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_replace))) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_do_read)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_do_read) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_valid_n <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_valid;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_first_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_first);
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_last_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_last);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_we <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_payload_we;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_addr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_sink_payload_addr;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_count <= 3'd4;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_ready <= 1'd1;
			end
		end
	end
	vns_bankmachine3_state <= vns_bankmachine3_next_state;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_close) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_opened <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_open) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_opened <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_replace))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_produce <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_do_read) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_consume <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_replace))) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_do_read)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_do_read) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_valid_n <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_valid;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_first_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_first);
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_last_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_last);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_we <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_payload_we;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_addr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_sink_payload_addr;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_count <= 3'd4;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_ready <= 1'd1;
			end
		end
	end
	vns_bankmachine4_state <= vns_bankmachine4_next_state;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_close) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_opened <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_open) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_opened <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_replace))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_produce <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_do_read) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_consume <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_replace))) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_do_read)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_do_read) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_valid_n <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_valid;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_first_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_first);
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_last_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_last);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_we <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_payload_we;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_addr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_sink_payload_addr;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_count <= 3'd4;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_ready <= 1'd1;
			end
		end
	end
	vns_bankmachine5_state <= vns_bankmachine5_next_state;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_close) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_opened <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_open) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_opened <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_replace))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_produce <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_do_read) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_consume <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_replace))) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_do_read)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_do_read) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_valid_n <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_valid;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_first_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_first);
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_last_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_last);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_we <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_payload_we;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_addr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_sink_payload_addr;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_count <= 3'd4;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_ready <= 1'd1;
			end
		end
	end
	vns_bankmachine6_state <= vns_bankmachine6_next_state;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_close) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_opened <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_open) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_opened <= 1'd1;
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_replace))) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_produce <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_do_read) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_consume <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_we & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable) & (~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_replace))) begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_do_read)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_do_read) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_level <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_valid_n <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_valid;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_first_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_first);
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_last_n <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_last);
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_pipe_ce) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_we <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_payload_we;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_addr <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_sink_payload_addr;
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_count <= 3'd5;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_count <= 3'd4;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_ready <= 1'd1;
			end
		end
	end
	vns_bankmachine7_state <= vns_bankmachine7_next_state;
	if ((~soc_videooverlaysoc_videooverlaysoc_sdram_en0)) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_time0 <= 5'd31;
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_max_time0)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_time0 <= (soc_videooverlaysoc_videooverlaysoc_sdram_time0 - 1'd1);
		end
	end
	if ((~soc_videooverlaysoc_videooverlaysoc_sdram_en1)) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_time1 <= 4'd15;
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_max_time1)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_time1 <= (soc_videooverlaysoc_videooverlaysoc_sdram_time1 - 1'd1);
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_ce) begin
		case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant)
			1'd0: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[1]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd1;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[2]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd2;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[3]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd3;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[4]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd4;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[5]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd5;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[6]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd6;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[7]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd7;
										end
									end
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[2]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd2;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[3]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd3;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[4]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd4;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[5]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd5;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[6]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd6;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[7]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd7;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[0]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd0;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[3]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd3;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[4]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd4;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[5]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd5;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[6]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd6;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[7]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd7;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[0]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd0;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[1]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd1;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[4]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd4;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[5]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd5;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[6]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd6;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[7]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd7;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[0]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd0;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[1]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd1;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[2]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd2;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[5]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd5;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[6]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd6;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[7]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd7;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[0]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd0;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[1]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd1;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[2]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd2;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[3]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd3;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[6]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd6;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[7]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd7;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[0]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd0;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[1]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd1;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[2]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd2;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[3]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd3;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[4]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd4;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd6: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[7]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd7;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[0]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd0;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[1]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd1;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[2]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd2;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[3]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd3;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[4]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd4;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[5]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd5;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd7: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[0]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd0;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[1]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 1'd1;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[2]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd2;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[3]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 2'd3;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[4]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd4;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[5]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd5;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_request[6]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd6;
										end
									end
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_ce) begin
		case (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant)
			1'd0: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[1]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd1;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[2]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd2;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[3]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd3;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[4]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd4;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[5]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd5;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[6]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd6;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[7]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd7;
										end
									end
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[2]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd2;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[3]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd3;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[4]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd4;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[5]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd5;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[6]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd6;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[7]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd7;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[0]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd0;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[3]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd3;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[4]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd4;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[5]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd5;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[6]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd6;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[7]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd7;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[0]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd0;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[1]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd1;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[4]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd4;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[5]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd5;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[6]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd6;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[7]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd7;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[0]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd0;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[1]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd1;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[2]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd2;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[5]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd5;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[6]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd6;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[7]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd7;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[0]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd0;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[1]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd1;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[2]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd2;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[3]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd3;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[6]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd6;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[7]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd7;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[0]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd0;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[1]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd1;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[2]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd2;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[3]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd3;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[4]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd4;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd6: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[7]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd7;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[0]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd0;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[1]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd1;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[2]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd2;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[3]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd3;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[4]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd4;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[5]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd5;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd7: begin
				if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[0]) begin
					soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd0;
				end else begin
					if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[1]) begin
						soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 1'd1;
					end else begin
						if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[2]) begin
							soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd2;
						end else begin
							if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[3]) begin
								soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 2'd3;
							end else begin
								if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[4]) begin
									soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd4;
								end else begin
									if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[5]) begin
										soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd5;
									end else begin
										if (soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_request[6]) begin
											soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd6;
										end
									end
								end
							end
						end
					end
				end
			end
		endcase
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cs_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_bank <= vns_sync_rhs_array_muxed0;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_address <= vns_sync_rhs_array_muxed1;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cas_n <= (~vns_sync_rhs_array_muxed2);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_ras_n <= (~vns_sync_rhs_array_muxed3);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_we_n <= (~vns_sync_rhs_array_muxed4);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_rddata_en <= vns_sync_rhs_array_muxed5;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_wrdata_en <= vns_sync_rhs_array_muxed6;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cs_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_bank <= vns_sync_rhs_array_muxed7;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_address <= vns_sync_rhs_array_muxed8;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cas_n <= (~vns_sync_rhs_array_muxed9);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_ras_n <= (~vns_sync_rhs_array_muxed10);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_we_n <= (~vns_sync_rhs_array_muxed11);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_rddata_en <= vns_sync_rhs_array_muxed12;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_wrdata_en <= vns_sync_rhs_array_muxed13;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cs_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_bank <= vns_sync_rhs_array_muxed14;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_address <= vns_sync_rhs_array_muxed15;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cas_n <= (~vns_sync_rhs_array_muxed16);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_ras_n <= (~vns_sync_rhs_array_muxed17);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_we_n <= (~vns_sync_rhs_array_muxed18);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_rddata_en <= vns_sync_rhs_array_muxed19;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_wrdata_en <= vns_sync_rhs_array_muxed20;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cs_n <= 1'd0;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_bank <= vns_sync_rhs_array_muxed21;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_address <= vns_sync_rhs_array_muxed22;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cas_n <= (~vns_sync_rhs_array_muxed23);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_ras_n <= (~vns_sync_rhs_array_muxed24);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_we_n <= (~vns_sync_rhs_array_muxed25);
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_rddata_en <= vns_sync_rhs_array_muxed26;
	soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_wrdata_en <= vns_sync_rhs_array_muxed27;
	if (soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_count <= 1'd1;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_ready <= 1'd1;
			end
		end
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_window <= {soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_window, soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_valid};
	if ((soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_count < 3'd4)) begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_count == 2'd3)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_ready <= (~soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_valid);
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_ready <= 1'd1;
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_count <= 1'd0;
		if (1'd1) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_ready <= 1'd1;
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_valid) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_count <= 3'd4;
		if (1'd0) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_ready <= 1'd1;
		end else begin
			soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_ready <= 1'd0;
		end
	end else begin
		if ((~soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_ready)) begin
			soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_count <= (soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_count - 1'd1);
			if ((soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_count == 1'd1)) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_ready <= 1'd1;
			end
		end
	end
	vns_multiplexer_state <= vns_multiplexer_next_state;
	soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_valid <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_valid;
	soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_ready <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_ready;
	soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_is_read <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_read;
	soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_is_write <= soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_cmd_payload_is_write;
	{soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_period, soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_counter} <= (soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_counter + 1'd1);
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_period) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads_r <= soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites_r <= soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites <= 1'd0;
	end else begin
		if ((soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_valid & soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_ready)) begin
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_is_read) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads <= (soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads + 1'd1);
			end
			if (soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_is_write) begin
				soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites <= (soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites + 1'd1);
			end
		end
	end
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_update_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads_status <= soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads_r;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites_status <= soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites_r;
	end
	if (((vns_roundrobin0_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_rdata_valid)) begin
		vns_rbank <= 1'd0;
	end
	if (((vns_roundrobin0_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_wdata_ready)) begin
		vns_wbank <= 1'd0;
	end
	if (((vns_roundrobin1_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_rdata_valid)) begin
		vns_rbank <= 1'd1;
	end
	if (((vns_roundrobin1_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_wdata_ready)) begin
		vns_wbank <= 1'd1;
	end
	if (((vns_roundrobin2_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_rdata_valid)) begin
		vns_rbank <= 2'd2;
	end
	if (((vns_roundrobin2_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_wdata_ready)) begin
		vns_wbank <= 2'd2;
	end
	if (((vns_roundrobin3_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_rdata_valid)) begin
		vns_rbank <= 2'd3;
	end
	if (((vns_roundrobin3_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_wdata_ready)) begin
		vns_wbank <= 2'd3;
	end
	if (((vns_roundrobin4_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_rdata_valid)) begin
		vns_rbank <= 3'd4;
	end
	if (((vns_roundrobin4_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_wdata_ready)) begin
		vns_wbank <= 3'd4;
	end
	if (((vns_roundrobin5_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_rdata_valid)) begin
		vns_rbank <= 3'd5;
	end
	if (((vns_roundrobin5_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_wdata_ready)) begin
		vns_wbank <= 3'd5;
	end
	if (((vns_roundrobin6_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_rdata_valid)) begin
		vns_rbank <= 3'd6;
	end
	if (((vns_roundrobin6_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_wdata_ready)) begin
		vns_wbank <= 3'd6;
	end
	if (((vns_roundrobin7_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_rdata_valid)) begin
		vns_rbank <= 3'd7;
	end
	if (((vns_roundrobin7_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_wdata_ready)) begin
		vns_wbank <= 3'd7;
	end
	vns_new_master_wdata_ready0 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_wdata_ready)) | ((vns_roundrobin1_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_wdata_ready)) | ((vns_roundrobin2_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_wdata_ready)) | ((vns_roundrobin3_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_wdata_ready)) | ((vns_roundrobin4_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_wdata_ready)) | ((vns_roundrobin5_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_wdata_ready)) | ((vns_roundrobin6_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_wdata_ready)) | ((vns_roundrobin7_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_wdata_ready));
	vns_new_master_wdata_ready1 <= vns_new_master_wdata_ready0;
	vns_new_master_wdata_ready2 <= vns_new_master_wdata_ready1;
	vns_new_master_wdata_ready3 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_wdata_ready)) | ((vns_roundrobin1_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_wdata_ready)) | ((vns_roundrobin2_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_wdata_ready)) | ((vns_roundrobin3_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_wdata_ready)) | ((vns_roundrobin4_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_wdata_ready)) | ((vns_roundrobin5_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_wdata_ready)) | ((vns_roundrobin6_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_wdata_ready)) | ((vns_roundrobin7_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_wdata_ready));
	vns_new_master_wdata_ready4 <= vns_new_master_wdata_ready3;
	vns_new_master_wdata_ready5 <= vns_new_master_wdata_ready4;
	vns_new_master_wdata_ready6 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_wdata_ready)) | ((vns_roundrobin1_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_wdata_ready)) | ((vns_roundrobin2_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_wdata_ready)) | ((vns_roundrobin3_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_wdata_ready)) | ((vns_roundrobin4_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_wdata_ready)) | ((vns_roundrobin5_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_wdata_ready)) | ((vns_roundrobin6_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_wdata_ready)) | ((vns_roundrobin7_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_wdata_ready));
	vns_new_master_wdata_ready7 <= vns_new_master_wdata_ready6;
	vns_new_master_wdata_ready8 <= vns_new_master_wdata_ready7;
	vns_new_master_rdata_valid0 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_rdata_valid)) | ((vns_roundrobin1_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_rdata_valid)) | ((vns_roundrobin2_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_rdata_valid)) | ((vns_roundrobin3_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_rdata_valid)) | ((vns_roundrobin4_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_rdata_valid)) | ((vns_roundrobin5_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_rdata_valid)) | ((vns_roundrobin6_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_rdata_valid)) | ((vns_roundrobin7_grant == 1'd0) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_rdata_valid));
	vns_new_master_rdata_valid1 <= vns_new_master_rdata_valid0;
	vns_new_master_rdata_valid2 <= vns_new_master_rdata_valid1;
	vns_new_master_rdata_valid3 <= vns_new_master_rdata_valid2;
	vns_new_master_rdata_valid4 <= vns_new_master_rdata_valid3;
	vns_new_master_rdata_valid5 <= vns_new_master_rdata_valid4;
	vns_new_master_rdata_valid6 <= vns_new_master_rdata_valid5;
	vns_new_master_rdata_valid7 <= vns_new_master_rdata_valid6;
	vns_new_master_rdata_valid8 <= vns_new_master_rdata_valid7;
	vns_new_master_rdata_valid9 <= vns_new_master_rdata_valid8;
	vns_new_master_rdata_valid10 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_rdata_valid)) | ((vns_roundrobin1_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_rdata_valid)) | ((vns_roundrobin2_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_rdata_valid)) | ((vns_roundrobin3_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_rdata_valid)) | ((vns_roundrobin4_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_rdata_valid)) | ((vns_roundrobin5_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_rdata_valid)) | ((vns_roundrobin6_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_rdata_valid)) | ((vns_roundrobin7_grant == 1'd1) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_rdata_valid));
	vns_new_master_rdata_valid11 <= vns_new_master_rdata_valid10;
	vns_new_master_rdata_valid12 <= vns_new_master_rdata_valid11;
	vns_new_master_rdata_valid13 <= vns_new_master_rdata_valid12;
	vns_new_master_rdata_valid14 <= vns_new_master_rdata_valid13;
	vns_new_master_rdata_valid15 <= vns_new_master_rdata_valid14;
	vns_new_master_rdata_valid16 <= vns_new_master_rdata_valid15;
	vns_new_master_rdata_valid17 <= vns_new_master_rdata_valid16;
	vns_new_master_rdata_valid18 <= vns_new_master_rdata_valid17;
	vns_new_master_rdata_valid19 <= vns_new_master_rdata_valid18;
	vns_new_master_rdata_valid20 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank0_rdata_valid)) | ((vns_roundrobin1_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank1_rdata_valid)) | ((vns_roundrobin2_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank2_rdata_valid)) | ((vns_roundrobin3_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank3_rdata_valid)) | ((vns_roundrobin4_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank4_rdata_valid)) | ((vns_roundrobin5_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank5_rdata_valid)) | ((vns_roundrobin6_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank6_rdata_valid)) | ((vns_roundrobin7_grant == 2'd2) & soc_videooverlaysoc_videooverlaysoc_sdram_interface_bank7_rdata_valid));
	vns_new_master_rdata_valid21 <= vns_new_master_rdata_valid20;
	vns_new_master_rdata_valid22 <= vns_new_master_rdata_valid21;
	vns_new_master_rdata_valid23 <= vns_new_master_rdata_valid22;
	vns_new_master_rdata_valid24 <= vns_new_master_rdata_valid23;
	vns_new_master_rdata_valid25 <= vns_new_master_rdata_valid24;
	vns_new_master_rdata_valid26 <= vns_new_master_rdata_valid25;
	vns_new_master_rdata_valid27 <= vns_new_master_rdata_valid26;
	vns_new_master_rdata_valid28 <= vns_new_master_rdata_valid27;
	vns_new_master_rdata_valid29 <= vns_new_master_rdata_valid28;
	soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_binary <= soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next_binary;
	soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q <= soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_next;
	soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_binary <= soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_next_binary;
	soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q <= soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_next;
	if (vns_roundrobin0_ce) begin
		case (vns_roundrobin0_grant)
			1'd0: begin
				if (vns_roundrobin0_request[1]) begin
					vns_roundrobin0_grant <= 1'd1;
				end else begin
					if (vns_roundrobin0_request[2]) begin
						vns_roundrobin0_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin0_request[2]) begin
					vns_roundrobin0_grant <= 2'd2;
				end else begin
					if (vns_roundrobin0_request[0]) begin
						vns_roundrobin0_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin0_request[0]) begin
					vns_roundrobin0_grant <= 1'd0;
				end else begin
					if (vns_roundrobin0_request[1]) begin
						vns_roundrobin0_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin1_ce) begin
		case (vns_roundrobin1_grant)
			1'd0: begin
				if (vns_roundrobin1_request[1]) begin
					vns_roundrobin1_grant <= 1'd1;
				end else begin
					if (vns_roundrobin1_request[2]) begin
						vns_roundrobin1_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin1_request[2]) begin
					vns_roundrobin1_grant <= 2'd2;
				end else begin
					if (vns_roundrobin1_request[0]) begin
						vns_roundrobin1_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin1_request[0]) begin
					vns_roundrobin1_grant <= 1'd0;
				end else begin
					if (vns_roundrobin1_request[1]) begin
						vns_roundrobin1_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin2_ce) begin
		case (vns_roundrobin2_grant)
			1'd0: begin
				if (vns_roundrobin2_request[1]) begin
					vns_roundrobin2_grant <= 1'd1;
				end else begin
					if (vns_roundrobin2_request[2]) begin
						vns_roundrobin2_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin2_request[2]) begin
					vns_roundrobin2_grant <= 2'd2;
				end else begin
					if (vns_roundrobin2_request[0]) begin
						vns_roundrobin2_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin2_request[0]) begin
					vns_roundrobin2_grant <= 1'd0;
				end else begin
					if (vns_roundrobin2_request[1]) begin
						vns_roundrobin2_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin3_ce) begin
		case (vns_roundrobin3_grant)
			1'd0: begin
				if (vns_roundrobin3_request[1]) begin
					vns_roundrobin3_grant <= 1'd1;
				end else begin
					if (vns_roundrobin3_request[2]) begin
						vns_roundrobin3_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin3_request[2]) begin
					vns_roundrobin3_grant <= 2'd2;
				end else begin
					if (vns_roundrobin3_request[0]) begin
						vns_roundrobin3_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin3_request[0]) begin
					vns_roundrobin3_grant <= 1'd0;
				end else begin
					if (vns_roundrobin3_request[1]) begin
						vns_roundrobin3_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin4_ce) begin
		case (vns_roundrobin4_grant)
			1'd0: begin
				if (vns_roundrobin4_request[1]) begin
					vns_roundrobin4_grant <= 1'd1;
				end else begin
					if (vns_roundrobin4_request[2]) begin
						vns_roundrobin4_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin4_request[2]) begin
					vns_roundrobin4_grant <= 2'd2;
				end else begin
					if (vns_roundrobin4_request[0]) begin
						vns_roundrobin4_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin4_request[0]) begin
					vns_roundrobin4_grant <= 1'd0;
				end else begin
					if (vns_roundrobin4_request[1]) begin
						vns_roundrobin4_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin5_ce) begin
		case (vns_roundrobin5_grant)
			1'd0: begin
				if (vns_roundrobin5_request[1]) begin
					vns_roundrobin5_grant <= 1'd1;
				end else begin
					if (vns_roundrobin5_request[2]) begin
						vns_roundrobin5_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin5_request[2]) begin
					vns_roundrobin5_grant <= 2'd2;
				end else begin
					if (vns_roundrobin5_request[0]) begin
						vns_roundrobin5_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin5_request[0]) begin
					vns_roundrobin5_grant <= 1'd0;
				end else begin
					if (vns_roundrobin5_request[1]) begin
						vns_roundrobin5_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin6_ce) begin
		case (vns_roundrobin6_grant)
			1'd0: begin
				if (vns_roundrobin6_request[1]) begin
					vns_roundrobin6_grant <= 1'd1;
				end else begin
					if (vns_roundrobin6_request[2]) begin
						vns_roundrobin6_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin6_request[2]) begin
					vns_roundrobin6_grant <= 2'd2;
				end else begin
					if (vns_roundrobin6_request[0]) begin
						vns_roundrobin6_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin6_request[0]) begin
					vns_roundrobin6_grant <= 1'd0;
				end else begin
					if (vns_roundrobin6_request[1]) begin
						vns_roundrobin6_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin7_ce) begin
		case (vns_roundrobin7_grant)
			1'd0: begin
				if (vns_roundrobin7_request[1]) begin
					vns_roundrobin7_grant <= 1'd1;
				end else begin
					if (vns_roundrobin7_request[2]) begin
						vns_roundrobin7_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin7_request[2]) begin
					vns_roundrobin7_grant <= 2'd2;
				end else begin
					if (vns_roundrobin7_request[0]) begin
						vns_roundrobin7_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin7_request[0]) begin
					vns_roundrobin7_grant <= 1'd0;
				end else begin
					if (vns_roundrobin7_request[1]) begin
						vns_roundrobin7_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	soc_videooverlaysoc_videooverlaysoc_adr_offset_r <= soc_videooverlaysoc_videooverlaysoc_interface0_wb_sdram_adr[2:0];
	vns_fullmemorywe_state <= vns_fullmemorywe_next_state;
	vns_litedramwishbone2native_state <= vns_litedramwishbone2native_next_state;
	if (soc_videooverlaysoc_hdmi_in0_freq_period_done) begin
		soc_videooverlaysoc_hdmi_in0_freq_period_counter <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in0_freq_period_counter <= (soc_videooverlaysoc_hdmi_in0_freq_period_counter + 1'd1);
	end
	soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o <= soc_videooverlaysoc_hdmi_in0_freq_gray_decoder_o_comb;
	soc_videooverlaysoc_hdmi_in0_freq_sampler_i_d <= soc_videooverlaysoc_hdmi_in0_freq_sampler_i;
	if (soc_videooverlaysoc_hdmi_in0_freq_sampler_latch) begin
		soc_videooverlaysoc_hdmi_in0_freq_sampler_counter <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_freq_sampler_o <= soc_videooverlaysoc_hdmi_in0_freq_sampler_counter;
	end else begin
		soc_videooverlaysoc_hdmi_in0_freq_sampler_counter <= (soc_videooverlaysoc_hdmi_in0_freq_sampler_counter + soc_videooverlaysoc_hdmi_in0_freq_sampler_inc);
	end
	soc_videooverlaysoc_hdmi_in0_edid_sda_drv_reg <= soc_videooverlaysoc_hdmi_in0_edid_sda_drv;
	{soc_videooverlaysoc_hdmi_in0_edid_samp_carry, soc_videooverlaysoc_hdmi_in0_edid_samp_count} <= (soc_videooverlaysoc_hdmi_in0_edid_samp_count + 1'd1);
	if (soc_videooverlaysoc_hdmi_in0_edid_samp_carry) begin
		soc_videooverlaysoc_hdmi_in0_edid_scl_i <= soc_videooverlaysoc_hdmi_in0_edid_scl_raw;
		soc_videooverlaysoc_hdmi_in0_edid_sda_i <= soc_videooverlaysoc_hdmi_in0_edid_sda_raw;
	end
	soc_videooverlaysoc_hdmi_in0_edid_scl_r <= soc_videooverlaysoc_hdmi_in0_edid_scl_i;
	soc_videooverlaysoc_hdmi_in0_edid_sda_r <= soc_videooverlaysoc_hdmi_in0_edid_sda_i;
	if (soc_videooverlaysoc_hdmi_in0_edid_start) begin
		soc_videooverlaysoc_hdmi_in0_edid_counter <= 1'd0;
	end
	if (soc_videooverlaysoc_hdmi_in0_edid_scl_rising) begin
		if ((soc_videooverlaysoc_hdmi_in0_edid_counter == 4'd8)) begin
			soc_videooverlaysoc_hdmi_in0_edid_counter <= 1'd0;
		end else begin
			soc_videooverlaysoc_hdmi_in0_edid_counter <= (soc_videooverlaysoc_hdmi_in0_edid_counter + 1'd1);
			soc_videooverlaysoc_hdmi_in0_edid_din <= {soc_videooverlaysoc_hdmi_in0_edid_din[6:0], soc_videooverlaysoc_hdmi_in0_edid_sda_i};
		end
	end
	if (soc_videooverlaysoc_hdmi_in0_edid_update_is_read) begin
		soc_videooverlaysoc_hdmi_in0_edid_is_read <= soc_videooverlaysoc_hdmi_in0_edid_din[0];
	end
	if (soc_videooverlaysoc_hdmi_in0_edid_oc_load) begin
		soc_videooverlaysoc_hdmi_in0_edid_offset_counter <= soc_videooverlaysoc_hdmi_in0_edid_din;
	end else begin
		if (soc_videooverlaysoc_hdmi_in0_edid_oc_inc) begin
			soc_videooverlaysoc_hdmi_in0_edid_offset_counter <= (soc_videooverlaysoc_hdmi_in0_edid_offset_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in0_edid_data_drv_en) begin
		soc_videooverlaysoc_hdmi_in0_edid_data_drv <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_hdmi_in0_edid_data_drv_stop) begin
			soc_videooverlaysoc_hdmi_in0_edid_data_drv <= 1'd0;
		end
	end
	if (soc_videooverlaysoc_hdmi_in0_edid_data_drv_en) begin
		case (soc_videooverlaysoc_hdmi_in0_edid_counter)
			1'd0: begin
				soc_videooverlaysoc_hdmi_in0_edid_data_bit <= soc_videooverlaysoc_hdmi_in0_edid_dat_r[7];
			end
			1'd1: begin
				soc_videooverlaysoc_hdmi_in0_edid_data_bit <= soc_videooverlaysoc_hdmi_in0_edid_dat_r[6];
			end
			2'd2: begin
				soc_videooverlaysoc_hdmi_in0_edid_data_bit <= soc_videooverlaysoc_hdmi_in0_edid_dat_r[5];
			end
			2'd3: begin
				soc_videooverlaysoc_hdmi_in0_edid_data_bit <= soc_videooverlaysoc_hdmi_in0_edid_dat_r[4];
			end
			3'd4: begin
				soc_videooverlaysoc_hdmi_in0_edid_data_bit <= soc_videooverlaysoc_hdmi_in0_edid_dat_r[3];
			end
			3'd5: begin
				soc_videooverlaysoc_hdmi_in0_edid_data_bit <= soc_videooverlaysoc_hdmi_in0_edid_dat_r[2];
			end
			3'd6: begin
				soc_videooverlaysoc_hdmi_in0_edid_data_bit <= soc_videooverlaysoc_hdmi_in0_edid_dat_r[1];
			end
			default: begin
				soc_videooverlaysoc_hdmi_in0_edid_data_bit <= soc_videooverlaysoc_hdmi_in0_edid_dat_r[0];
			end
		endcase
	end
	vns_edid0_state <= vns_edid0_next_state;
	if ((soc_videooverlaysoc_hdmi_in0_mmcm_read_re | soc_videooverlaysoc_hdmi_in0_mmcm_write_re)) begin
		soc_videooverlaysoc_hdmi_in0_mmcm_drdy_status <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in0_mmcm_drdy) begin
			soc_videooverlaysoc_hdmi_in0_mmcm_drdy_status <= 1'd1;
		end
	end
	if ((soc_videooverlaysoc_hdmi_in0_mmcm_read_o_re | soc_videooverlaysoc_hdmi_in0_mmcm_write_o_re)) begin
		soc_videooverlaysoc_hdmi_in0_mmcm_drdy_o_status <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in0_mmcm_drdy_o) begin
			soc_videooverlaysoc_hdmi_in0_mmcm_drdy_o_status <= 1'd1;
		end
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_rst_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_master_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_delay_slave_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture0_do_reset_lateness_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_wer0_o) begin
		soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_sys <= soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_r;
	end
	if (soc_videooverlaysoc_hdmi_in0_wer0_update_re) begin
		soc_videooverlaysoc_hdmi_in0_wer0_status <= soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_sys;
	end
	soc_videooverlaysoc_hdmi_in0_wer0_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_wer0_toggle_o;
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_rst_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_master_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_delay_slave_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture1_do_reset_lateness_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_wer1_o) begin
		soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_sys <= soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_r;
	end
	if (soc_videooverlaysoc_hdmi_in0_wer1_update_re) begin
		soc_videooverlaysoc_hdmi_in0_wer1_status <= soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_sys;
	end
	soc_videooverlaysoc_hdmi_in0_wer1_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_wer1_toggle_o;
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_rst_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_master_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_delay_slave_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_i) begin
		soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_i <= (~soc_videooverlaysoc_hdmi_in0_s7datacapture2_do_reset_lateness_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in0_wer2_o) begin
		soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_sys <= soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_r;
	end
	if (soc_videooverlaysoc_hdmi_in0_wer2_update_re) begin
		soc_videooverlaysoc_hdmi_in0_wer2_status <= soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_sys;
	end
	soc_videooverlaysoc_hdmi_in0_wer2_toggle_o_r <= soc_videooverlaysoc_hdmi_in0_wer2_toggle_o;
	if (soc_videooverlaysoc_hdmi_in1_freq_period_done) begin
		soc_videooverlaysoc_hdmi_in1_freq_period_counter <= 1'd0;
	end else begin
		soc_videooverlaysoc_hdmi_in1_freq_period_counter <= (soc_videooverlaysoc_hdmi_in1_freq_period_counter + 1'd1);
	end
	soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o <= soc_videooverlaysoc_hdmi_in1_freq_gray_decoder_o_comb;
	soc_videooverlaysoc_hdmi_in1_freq_sampler_i_d <= soc_videooverlaysoc_hdmi_in1_freq_sampler_i;
	if (soc_videooverlaysoc_hdmi_in1_freq_sampler_latch) begin
		soc_videooverlaysoc_hdmi_in1_freq_sampler_counter <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_freq_sampler_o <= soc_videooverlaysoc_hdmi_in1_freq_sampler_counter;
	end else begin
		soc_videooverlaysoc_hdmi_in1_freq_sampler_counter <= (soc_videooverlaysoc_hdmi_in1_freq_sampler_counter + soc_videooverlaysoc_hdmi_in1_freq_sampler_inc);
	end
	soc_videooverlaysoc_hdmi_in1_edid_sda_drv_reg <= soc_videooverlaysoc_hdmi_in1_edid_sda_drv;
	{soc_videooverlaysoc_hdmi_in1_edid_samp_carry, soc_videooverlaysoc_hdmi_in1_edid_samp_count} <= (soc_videooverlaysoc_hdmi_in1_edid_samp_count + 1'd1);
	if (soc_videooverlaysoc_hdmi_in1_edid_samp_carry) begin
		soc_videooverlaysoc_hdmi_in1_edid_scl_i <= soc_videooverlaysoc_hdmi_in1_edid_scl_raw;
		soc_videooverlaysoc_hdmi_in1_edid_sda_i <= soc_videooverlaysoc_hdmi_in1_edid_sda_raw;
	end
	soc_videooverlaysoc_hdmi_in1_edid_scl_r <= soc_videooverlaysoc_hdmi_in1_edid_scl_i;
	soc_videooverlaysoc_hdmi_in1_edid_sda_r <= soc_videooverlaysoc_hdmi_in1_edid_sda_i;
	if (soc_videooverlaysoc_hdmi_in1_edid_start) begin
		soc_videooverlaysoc_hdmi_in1_edid_counter <= 1'd0;
	end
	if (soc_videooverlaysoc_hdmi_in1_edid_scl_rising) begin
		if ((soc_videooverlaysoc_hdmi_in1_edid_counter == 4'd8)) begin
			soc_videooverlaysoc_hdmi_in1_edid_counter <= 1'd0;
		end else begin
			soc_videooverlaysoc_hdmi_in1_edid_counter <= (soc_videooverlaysoc_hdmi_in1_edid_counter + 1'd1);
			soc_videooverlaysoc_hdmi_in1_edid_din <= {soc_videooverlaysoc_hdmi_in1_edid_din[6:0], soc_videooverlaysoc_hdmi_in1_edid_sda_i};
		end
	end
	if (soc_videooverlaysoc_hdmi_in1_edid_update_is_read) begin
		soc_videooverlaysoc_hdmi_in1_edid_is_read <= soc_videooverlaysoc_hdmi_in1_edid_din[0];
	end
	if (soc_videooverlaysoc_hdmi_in1_edid_oc_load) begin
		soc_videooverlaysoc_hdmi_in1_edid_offset_counter <= soc_videooverlaysoc_hdmi_in1_edid_din;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_edid_oc_inc) begin
			soc_videooverlaysoc_hdmi_in1_edid_offset_counter <= (soc_videooverlaysoc_hdmi_in1_edid_offset_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in1_edid_data_drv_en) begin
		soc_videooverlaysoc_hdmi_in1_edid_data_drv <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_edid_data_drv_stop) begin
			soc_videooverlaysoc_hdmi_in1_edid_data_drv <= 1'd0;
		end
	end
	if (soc_videooverlaysoc_hdmi_in1_edid_data_drv_en) begin
		case (soc_videooverlaysoc_hdmi_in1_edid_counter)
			1'd0: begin
				soc_videooverlaysoc_hdmi_in1_edid_data_bit <= soc_videooverlaysoc_hdmi_in1_edid_dat_r[7];
			end
			1'd1: begin
				soc_videooverlaysoc_hdmi_in1_edid_data_bit <= soc_videooverlaysoc_hdmi_in1_edid_dat_r[6];
			end
			2'd2: begin
				soc_videooverlaysoc_hdmi_in1_edid_data_bit <= soc_videooverlaysoc_hdmi_in1_edid_dat_r[5];
			end
			2'd3: begin
				soc_videooverlaysoc_hdmi_in1_edid_data_bit <= soc_videooverlaysoc_hdmi_in1_edid_dat_r[4];
			end
			3'd4: begin
				soc_videooverlaysoc_hdmi_in1_edid_data_bit <= soc_videooverlaysoc_hdmi_in1_edid_dat_r[3];
			end
			3'd5: begin
				soc_videooverlaysoc_hdmi_in1_edid_data_bit <= soc_videooverlaysoc_hdmi_in1_edid_dat_r[2];
			end
			3'd6: begin
				soc_videooverlaysoc_hdmi_in1_edid_data_bit <= soc_videooverlaysoc_hdmi_in1_edid_dat_r[1];
			end
			default: begin
				soc_videooverlaysoc_hdmi_in1_edid_data_bit <= soc_videooverlaysoc_hdmi_in1_edid_dat_r[0];
			end
		endcase
	end
	vns_edid1_state <= vns_edid1_next_state;
	if ((soc_videooverlaysoc_hdmi_in1_mmcm_read_re | soc_videooverlaysoc_hdmi_in1_mmcm_write_re)) begin
		soc_videooverlaysoc_hdmi_in1_mmcm_drdy_status <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_mmcm_drdy) begin
			soc_videooverlaysoc_hdmi_in1_mmcm_drdy_status <= 1'd1;
		end
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_rst_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_master_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_delay_slave_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture0_do_reset_lateness_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_wer0_o) begin
		soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_sys <= soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_r;
	end
	if (soc_videooverlaysoc_hdmi_in1_wer0_update_re) begin
		soc_videooverlaysoc_hdmi_in1_wer0_status <= soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_sys;
	end
	soc_videooverlaysoc_hdmi_in1_wer0_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_wer0_toggle_o;
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_rst_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_master_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_delay_slave_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture1_do_reset_lateness_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_wer1_o) begin
		soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_sys <= soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_r;
	end
	if (soc_videooverlaysoc_hdmi_in1_wer1_update_re) begin
		soc_videooverlaysoc_hdmi_in1_wer1_status <= soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_sys;
	end
	soc_videooverlaysoc_hdmi_in1_wer1_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_wer1_toggle_o;
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_rst_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_master_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_inc_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_delay_slave_dec_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_i) begin
		soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_s7datacapture2_do_reset_lateness_toggle_i);
	end
	if (soc_videooverlaysoc_hdmi_in1_wer2_o) begin
		soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_sys <= soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_r;
	end
	if (soc_videooverlaysoc_hdmi_in1_wer2_update_re) begin
		soc_videooverlaysoc_hdmi_in1_wer2_status <= soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_sys;
	end
	soc_videooverlaysoc_hdmi_in1_wer2_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_wer2_toggle_o;
	if (soc_videooverlaysoc_hdmi_in1_frame_overflow_re) begin
		soc_videooverlaysoc_hdmi_in1_frame_overflow_mask <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_o) begin
			soc_videooverlaysoc_hdmi_in1_frame_overflow_mask <= 1'd0;
		end
	end
	soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_binary <= soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next_binary;
	soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q <= soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_next;
	if (soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_i) begin
		soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_i <= (~soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_toggle_i);
	end
	soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_o_r <= soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_o;
	if (soc_videooverlaysoc_hdmi_in1_dma_reset_words) begin
		soc_videooverlaysoc_hdmi_in1_dma_current_address <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_address;
		soc_videooverlaysoc_hdmi_in1_dma_mwords_remaining <= soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage;
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_dma_count_word) begin
			soc_videooverlaysoc_hdmi_in1_dma_current_address <= (soc_videooverlaysoc_hdmi_in1_dma_current_address + 1'd1);
			soc_videooverlaysoc_hdmi_in1_dma_mwords_remaining <= (soc_videooverlaysoc_hdmi_in1_dma_mwords_remaining - 1'd1);
		end
	end
	if (soc_videooverlaysoc_hdmi_in1_dma_slot_array_change_slot) begin
		if (soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_valid) begin
			soc_videooverlaysoc_hdmi_in1_dma_slot_array_current_slot <= 1'd1;
		end
		if (soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_valid) begin
			soc_videooverlaysoc_hdmi_in1_dma_slot_array_current_slot <= 1'd0;
		end
	end
	if (((soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_we & soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_writable) & (~soc_videooverlaysoc_hdmi_in1_dma_fifo_replace))) begin
		soc_videooverlaysoc_hdmi_in1_dma_fifo_produce <= (soc_videooverlaysoc_hdmi_in1_dma_fifo_produce + 1'd1);
	end
	if (soc_videooverlaysoc_hdmi_in1_dma_fifo_do_read) begin
		soc_videooverlaysoc_hdmi_in1_dma_fifo_consume <= (soc_videooverlaysoc_hdmi_in1_dma_fifo_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_we & soc_videooverlaysoc_hdmi_in1_dma_fifo_syncfifo_writable) & (~soc_videooverlaysoc_hdmi_in1_dma_fifo_replace))) begin
		if ((~soc_videooverlaysoc_hdmi_in1_dma_fifo_do_read)) begin
			soc_videooverlaysoc_hdmi_in1_dma_fifo_level <= (soc_videooverlaysoc_hdmi_in1_dma_fifo_level + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_hdmi_in1_dma_fifo_do_read) begin
			soc_videooverlaysoc_hdmi_in1_dma_fifo_level <= (soc_videooverlaysoc_hdmi_in1_dma_fifo_level - 1'd1);
		end
	end
	vns_dma_state <= vns_dma_next_state;
	soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_binary <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_next_binary;
	soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_next;
	if (soc_videooverlaysoc_hdmi_core_out0_i) begin
		soc_videooverlaysoc_hdmi_core_out0_toggle_i <= (~soc_videooverlaysoc_hdmi_core_out0_toggle_i);
	end
	if (soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter_reset) begin
		soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter_ce) begin
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter <= (soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_load) begin
		soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header_reg <= soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header;
	end else begin
		if (soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_shift) begin
			soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header_reg <= {soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer, soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_header_reg[63:32]};
		end
	end
	vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_state <= vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_next_state;
	vns_liteethetherbonepackettx_fsm_state <= vns_liteethetherbonepackettx_fsm_next_state;
	soc_videooverlaysoc_packet_valid <= (soc_videooverlaysoc_packet_depacketizer_source_valid & (soc_videooverlaysoc_packet_depacketizer_source_param_magic == 15'd20079));
	if (soc_videooverlaysoc_packet_depacketizer_counter_reset) begin
		soc_videooverlaysoc_packet_depacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_packet_depacketizer_counter_ce) begin
			soc_videooverlaysoc_packet_depacketizer_counter <= (soc_videooverlaysoc_packet_depacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_packet_depacketizer_shift) begin
		soc_videooverlaysoc_packet_depacketizer_header_reg <= {soc_videooverlaysoc_packet_depacketizer_sink_payload_data, soc_videooverlaysoc_packet_depacketizer_header_reg[63:32]};
	end
	if (soc_videooverlaysoc_packet_depacketizer_is_el) begin
		soc_videooverlaysoc_packet_depacketizer_no_payload <= soc_videooverlaysoc_packet_depacketizer_sink_last;
	end
	vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_state <= vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_next_state;
	vns_liteethetherbonepacketrx_fsm_state <= vns_liteethetherbonepacketrx_fsm_next_state;
	vns_liteethetherboneprobe_state <= vns_liteethetherboneprobe_next_state;
	if ((soc_videooverlaysoc_record_sink_sink_valid & soc_videooverlaysoc_record_sink_sink_ready)) begin
		if (soc_videooverlaysoc_record_first) begin
			soc_videooverlaysoc_record_last_ip_address <= soc_videooverlaysoc_record_sink_sink_param_ip_address;
		end
		soc_videooverlaysoc_record_first <= soc_videooverlaysoc_record_sink_sink_last;
	end
	if (soc_videooverlaysoc_record_depacketizer_counter_reset) begin
		soc_videooverlaysoc_record_depacketizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_record_depacketizer_counter_ce) begin
			soc_videooverlaysoc_record_depacketizer_counter <= (soc_videooverlaysoc_record_depacketizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_record_depacketizer_shift) begin
		soc_videooverlaysoc_record_depacketizer_header_reg <= soc_videooverlaysoc_record_depacketizer_sink_payload_data;
	end
	if (soc_videooverlaysoc_record_depacketizer_is_el) begin
		soc_videooverlaysoc_record_depacketizer_no_payload <= soc_videooverlaysoc_record_depacketizer_sink_last;
	end
	vns_liteethetherbonerecorddepacketizer_state <= vns_liteethetherbonerecorddepacketizer_next_state;
	if (soc_videooverlaysoc_record_receiver_base_addr_update) begin
		soc_videooverlaysoc_record_receiver_base_addr <= soc_videooverlaysoc_record_receiver_fifo_source_payload_data;
	end
	if (soc_videooverlaysoc_record_receiver_counter_reset) begin
		soc_videooverlaysoc_record_receiver_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_record_receiver_counter_ce) begin
			soc_videooverlaysoc_record_receiver_counter <= (soc_videooverlaysoc_record_receiver_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_record_receiver_fifo_syncfifo_re) begin
		soc_videooverlaysoc_record_receiver_fifo_readable <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_record_receiver_fifo_re) begin
			soc_videooverlaysoc_record_receiver_fifo_readable <= 1'd0;
		end
	end
	if (((soc_videooverlaysoc_record_receiver_fifo_syncfifo_we & soc_videooverlaysoc_record_receiver_fifo_syncfifo_writable) & (~soc_videooverlaysoc_record_receiver_fifo_replace))) begin
		soc_videooverlaysoc_record_receiver_fifo_produce <= (soc_videooverlaysoc_record_receiver_fifo_produce + 1'd1);
	end
	if (soc_videooverlaysoc_record_receiver_fifo_do_read) begin
		soc_videooverlaysoc_record_receiver_fifo_consume <= (soc_videooverlaysoc_record_receiver_fifo_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_record_receiver_fifo_syncfifo_we & soc_videooverlaysoc_record_receiver_fifo_syncfifo_writable) & (~soc_videooverlaysoc_record_receiver_fifo_replace))) begin
		if ((~soc_videooverlaysoc_record_receiver_fifo_do_read)) begin
			soc_videooverlaysoc_record_receiver_fifo_level0 <= (soc_videooverlaysoc_record_receiver_fifo_level0 + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_record_receiver_fifo_do_read) begin
			soc_videooverlaysoc_record_receiver_fifo_level0 <= (soc_videooverlaysoc_record_receiver_fifo_level0 - 1'd1);
		end
	end
	vns_liteethetherbonerecordreceiver_state <= vns_liteethetherbonerecordreceiver_next_state;
	soc_videooverlaysoc_record_sender_source_source_param_byte_enable <= soc_videooverlaysoc_record_sender_fifo_source_param_be;
	if (soc_videooverlaysoc_record_sender_fifo_source_param_we) begin
		soc_videooverlaysoc_record_sender_source_source_param_wcount <= soc_videooverlaysoc_record_sender_fifo_source_param_count;
	end else begin
		soc_videooverlaysoc_record_sender_source_source_param_rcount <= soc_videooverlaysoc_record_sender_fifo_source_param_count;
	end
	if (soc_videooverlaysoc_record_sender_data_sel) begin
		soc_videooverlaysoc_record_sender_source_source_payload_data <= soc_videooverlaysoc_record_sender_fifo_source_payload_data;
	end else begin
		soc_videooverlaysoc_record_sender_source_source_payload_data <= soc_videooverlaysoc_record_sender_fifo_source_param_base_addr;
	end
	if (soc_videooverlaysoc_record_sender_fifo_syncfifo_re) begin
		soc_videooverlaysoc_record_sender_fifo_readable <= 1'd1;
	end else begin
		if (soc_videooverlaysoc_record_sender_fifo_re) begin
			soc_videooverlaysoc_record_sender_fifo_readable <= 1'd0;
		end
	end
	if (((soc_videooverlaysoc_record_sender_fifo_syncfifo_we & soc_videooverlaysoc_record_sender_fifo_syncfifo_writable) & (~soc_videooverlaysoc_record_sender_fifo_replace))) begin
		soc_videooverlaysoc_record_sender_fifo_produce <= (soc_videooverlaysoc_record_sender_fifo_produce + 1'd1);
	end
	if (soc_videooverlaysoc_record_sender_fifo_do_read) begin
		soc_videooverlaysoc_record_sender_fifo_consume <= (soc_videooverlaysoc_record_sender_fifo_consume + 1'd1);
	end
	if (((soc_videooverlaysoc_record_sender_fifo_syncfifo_we & soc_videooverlaysoc_record_sender_fifo_syncfifo_writable) & (~soc_videooverlaysoc_record_sender_fifo_replace))) begin
		if ((~soc_videooverlaysoc_record_sender_fifo_do_read)) begin
			soc_videooverlaysoc_record_sender_fifo_level0 <= (soc_videooverlaysoc_record_sender_fifo_level0 + 1'd1);
		end
	end else begin
		if (soc_videooverlaysoc_record_sender_fifo_do_read) begin
			soc_videooverlaysoc_record_sender_fifo_level0 <= (soc_videooverlaysoc_record_sender_fifo_level0 - 1'd1);
		end
	end
	vns_liteethetherbonerecordsender_state <= vns_liteethetherbonerecordsender_next_state;
	if (soc_videooverlaysoc_record_packetizer_counter_reset) begin
		soc_videooverlaysoc_record_packetizer_counter <= 1'd0;
	end else begin
		if (soc_videooverlaysoc_record_packetizer_counter_ce) begin
			soc_videooverlaysoc_record_packetizer_counter <= (soc_videooverlaysoc_record_packetizer_counter + 1'd1);
		end
	end
	if (soc_videooverlaysoc_record_packetizer_load) begin
		soc_videooverlaysoc_record_packetizer_header_reg <= soc_videooverlaysoc_record_packetizer_header;
	end
	vns_liteethetherbonerecordpacketizer_state <= vns_liteethetherbonerecordpacketizer_next_state;
	if (soc_videooverlaysoc_dispatcher_first) begin
		soc_videooverlaysoc_dispatcher_sel_ongoing <= soc_videooverlaysoc_dispatcher_sel0;
	end
	soc_videooverlaysoc_dispatcher_ongoing1 <= ((soc_videooverlaysoc_packet_source_source_valid | soc_videooverlaysoc_dispatcher_ongoing1) & (~soc_videooverlaysoc_dispatcher_last));
	if (soc_videooverlaysoc_dispatcher_last) begin
		soc_videooverlaysoc_dispatcher_first <= 1'd1;
	end else begin
		if ((soc_videooverlaysoc_packet_source_source_valid & soc_videooverlaysoc_packet_source_source_ready)) begin
			soc_videooverlaysoc_dispatcher_first <= 1'd0;
		end
	end
	case (soc_videooverlaysoc_grant)
		1'd0: begin
			if ((~soc_videooverlaysoc_request[0])) begin
				if (soc_videooverlaysoc_request[1]) begin
					soc_videooverlaysoc_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~soc_videooverlaysoc_request[1])) begin
				if (soc_videooverlaysoc_request[0]) begin
					soc_videooverlaysoc_grant <= 1'd0;
				end
			end
		end
	endcase
	soc_videooverlaysoc_status0_ongoing1 <= ((soc_videooverlaysoc_probe_source_valid | soc_videooverlaysoc_status0_ongoing1) & (~soc_videooverlaysoc_status0_last));
	if (soc_videooverlaysoc_status0_last) begin
		soc_videooverlaysoc_status0_first <= 1'd1;
	end else begin
		if ((soc_videooverlaysoc_probe_source_valid & soc_videooverlaysoc_probe_source_ready)) begin
			soc_videooverlaysoc_status0_first <= 1'd0;
		end
	end
	soc_videooverlaysoc_status1_ongoing1 <= ((soc_videooverlaysoc_record_source_source_valid | soc_videooverlaysoc_status1_ongoing1) & (~soc_videooverlaysoc_status1_last));
	if (soc_videooverlaysoc_status1_last) begin
		soc_videooverlaysoc_status1_first <= 1'd1;
	end else begin
		if ((soc_videooverlaysoc_record_source_source_valid & soc_videooverlaysoc_record_source_source_ready)) begin
			soc_videooverlaysoc_status1_first <= 1'd0;
		end
	end
	soc_videooverlaysoc_wishbone_source_param_base_addr <= soc_videooverlaysoc_wishbone_sink_param_base_addr;
	soc_videooverlaysoc_wishbone_source_payload_addr <= soc_videooverlaysoc_wishbone_sink_payload_addr;
	soc_videooverlaysoc_wishbone_source_param_count <= soc_videooverlaysoc_wishbone_sink_param_count;
	soc_videooverlaysoc_wishbone_source_param_be <= soc_videooverlaysoc_wishbone_sink_param_be;
	soc_videooverlaysoc_wishbone_source_param_we <= 1'd1;
	if (soc_videooverlaysoc_wishbone_data_update) begin
		soc_videooverlaysoc_wishbone_source_payload_data <= soc_videooverlaysoc_wishbone_bus_dat_r;
	end
	vns_liteethetherbonewishbonemaster_state <= vns_liteethetherbonewishbonemaster_next_state;
	case (vns_videooverlaysoc_grant)
		1'd0: begin
			if ((~vns_videooverlaysoc_request[0])) begin
				if (vns_videooverlaysoc_request[1]) begin
					vns_videooverlaysoc_grant <= 1'd1;
				end else begin
					if (vns_videooverlaysoc_request[2]) begin
						vns_videooverlaysoc_grant <= 2'd2;
					end
				end
			end
		end
		1'd1: begin
			if ((~vns_videooverlaysoc_request[1])) begin
				if (vns_videooverlaysoc_request[2]) begin
					vns_videooverlaysoc_grant <= 2'd2;
				end else begin
					if (vns_videooverlaysoc_request[0]) begin
						vns_videooverlaysoc_grant <= 1'd0;
					end
				end
			end
		end
		2'd2: begin
			if ((~vns_videooverlaysoc_request[2])) begin
				if (vns_videooverlaysoc_request[0]) begin
					vns_videooverlaysoc_grant <= 1'd0;
				end else begin
					if (vns_videooverlaysoc_request[1]) begin
						vns_videooverlaysoc_grant <= 1'd1;
					end
				end
			end
		end
	endcase
	vns_videooverlaysoc_slave_sel_r <= vns_videooverlaysoc_slave_sel;
	if (vns_videooverlaysoc_wait) begin
		if ((~vns_videooverlaysoc_done)) begin
			vns_videooverlaysoc_count <= (vns_videooverlaysoc_count - 1'd1);
		end
	end else begin
		vns_videooverlaysoc_count <= 17'd65536;
	end
	vns_videooverlaysoc_interface0_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank0_sel) begin
		case (vns_videooverlaysoc_interface0_bank_bus_adr[3:0])
			1'd0: begin
				vns_videooverlaysoc_interface0_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_reset_reset_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface0_bank_bus_dat_r <= vns_videooverlaysoc_csrbank0_scratch3_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface0_bank_bus_dat_r <= vns_videooverlaysoc_csrbank0_scratch2_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface0_bank_bus_dat_r <= vns_videooverlaysoc_csrbank0_scratch1_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface0_bank_bus_dat_r <= vns_videooverlaysoc_csrbank0_scratch0_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface0_bank_bus_dat_r <= vns_videooverlaysoc_csrbank0_bus_errors3_w;
			end
			3'd6: begin
				vns_videooverlaysoc_interface0_bank_bus_dat_r <= vns_videooverlaysoc_csrbank0_bus_errors2_w;
			end
			3'd7: begin
				vns_videooverlaysoc_interface0_bank_bus_dat_r <= vns_videooverlaysoc_csrbank0_bus_errors1_w;
			end
			4'd8: begin
				vns_videooverlaysoc_interface0_bank_bus_dat_r <= vns_videooverlaysoc_csrbank0_bus_errors0_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank0_scratch3_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full[31:24] <= vns_videooverlaysoc_csrbank0_scratch3_r;
	end
	if (vns_videooverlaysoc_csrbank0_scratch2_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full[23:16] <= vns_videooverlaysoc_csrbank0_scratch2_r;
	end
	if (vns_videooverlaysoc_csrbank0_scratch1_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full[15:8] <= vns_videooverlaysoc_csrbank0_scratch1_r;
	end
	if (vns_videooverlaysoc_csrbank0_scratch0_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full[7:0] <= vns_videooverlaysoc_csrbank0_scratch0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_re <= vns_videooverlaysoc_csrbank0_scratch0_re;
	vns_videooverlaysoc_interface1_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank1_sel) begin
		case (vns_videooverlaysoc_interface1_bank_bus_adr[2:0])
			1'd0: begin
				vns_videooverlaysoc_interface1_bank_bus_dat_r <= vns_videooverlaysoc_csrbank1_half_sys8x_taps0_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface1_bank_bus_dat_r <= vns_videooverlaysoc_csrbank1_dly_sel0_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface1_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface1_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface1_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_rst_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface1_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_bitslip_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank1_half_sys8x_taps0_re) begin
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_half_sys8x_taps_storage_full[3:0] <= vns_videooverlaysoc_csrbank1_half_sys8x_taps0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_half_sys8x_taps_re <= vns_videooverlaysoc_csrbank1_half_sys8x_taps0_re;
	if (vns_videooverlaysoc_csrbank1_dly_sel0_re) begin
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage_full[3:0] <= vns_videooverlaysoc_csrbank1_dly_sel0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_re <= vns_videooverlaysoc_csrbank1_dly_sel0_re;
	vns_videooverlaysoc_interface2_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank2_sel) begin
		case (vns_videooverlaysoc_interface2_bank_bus_adr[3:0])
			1'd0: begin
				vns_videooverlaysoc_interface2_bank_bus_dat_r <= vns_videooverlaysoc_csrbank2_Km6_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface2_bank_bus_dat_r <= vns_videooverlaysoc_csrbank2_Km5_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface2_bank_bus_dat_r <= vns_videooverlaysoc_csrbank2_Km4_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface2_bank_bus_dat_r <= vns_videooverlaysoc_csrbank2_Km3_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface2_bank_bus_dat_r <= vns_videooverlaysoc_csrbank2_Km2_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface2_bank_bus_dat_r <= vns_videooverlaysoc_csrbank2_Km1_w;
			end
			3'd6: begin
				vns_videooverlaysoc_interface2_bank_bus_dat_r <= vns_videooverlaysoc_csrbank2_Km0_w;
			end
			3'd7: begin
				vns_videooverlaysoc_interface2_bank_bus_dat_r <= vns_videooverlaysoc_csrbank2_Km_valid0_w;
			end
			4'd8: begin
				vns_videooverlaysoc_interface2_bank_bus_dat_r <= vns_videooverlaysoc_csrbank2_hpd_ena0_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank2_Km6_re) begin
		soc_videooverlaysoc_hdcp_Km_storage_full[55:48] <= vns_videooverlaysoc_csrbank2_Km6_r;
	end
	if (vns_videooverlaysoc_csrbank2_Km5_re) begin
		soc_videooverlaysoc_hdcp_Km_storage_full[47:40] <= vns_videooverlaysoc_csrbank2_Km5_r;
	end
	if (vns_videooverlaysoc_csrbank2_Km4_re) begin
		soc_videooverlaysoc_hdcp_Km_storage_full[39:32] <= vns_videooverlaysoc_csrbank2_Km4_r;
	end
	if (vns_videooverlaysoc_csrbank2_Km3_re) begin
		soc_videooverlaysoc_hdcp_Km_storage_full[31:24] <= vns_videooverlaysoc_csrbank2_Km3_r;
	end
	if (vns_videooverlaysoc_csrbank2_Km2_re) begin
		soc_videooverlaysoc_hdcp_Km_storage_full[23:16] <= vns_videooverlaysoc_csrbank2_Km2_r;
	end
	if (vns_videooverlaysoc_csrbank2_Km1_re) begin
		soc_videooverlaysoc_hdcp_Km_storage_full[15:8] <= vns_videooverlaysoc_csrbank2_Km1_r;
	end
	if (vns_videooverlaysoc_csrbank2_Km0_re) begin
		soc_videooverlaysoc_hdcp_Km_storage_full[7:0] <= vns_videooverlaysoc_csrbank2_Km0_r;
	end
	soc_videooverlaysoc_hdcp_Km_re <= vns_videooverlaysoc_csrbank2_Km0_re;
	if (vns_videooverlaysoc_csrbank2_Km_valid0_re) begin
		soc_videooverlaysoc_hdcp_Km_valid_storage_full <= vns_videooverlaysoc_csrbank2_Km_valid0_r;
	end
	soc_videooverlaysoc_hdcp_Km_valid_re <= vns_videooverlaysoc_csrbank2_Km_valid0_re;
	if (vns_videooverlaysoc_csrbank2_hpd_ena0_re) begin
		soc_videooverlaysoc_hdcp_hpd_ena_storage_full <= vns_videooverlaysoc_csrbank2_hpd_ena0_r;
	end
	soc_videooverlaysoc_hdcp_hpd_ena_re <= vns_videooverlaysoc_csrbank2_hpd_ena0_re;
	vns_videooverlaysoc_interface3_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank3_sel) begin
		case (vns_videooverlaysoc_interface3_bank_bus_adr[5:0])
			1'd0: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_underflow_enable0_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_core_out0_underflow_update_underflow_update_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_underflow_counter3_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_underflow_counter2_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_underflow_counter1_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_underflow_counter0_w;
			end
			3'd6: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_enable0_w;
			end
			3'd7: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_hres1_w;
			end
			4'd8: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_hres0_w;
			end
			4'd9: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_hsync_start1_w;
			end
			4'd10: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_hsync_start0_w;
			end
			4'd11: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_hsync_end1_w;
			end
			4'd12: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_hsync_end0_w;
			end
			4'd13: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_hscan1_w;
			end
			4'd14: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_hscan0_w;
			end
			4'd15: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_vres1_w;
			end
			5'd16: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_vres0_w;
			end
			5'd17: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_vsync_start1_w;
			end
			5'd18: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_vsync_start0_w;
			end
			5'd19: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_vsync_end1_w;
			end
			5'd20: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_vsync_end0_w;
			end
			5'd21: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_vscan1_w;
			end
			5'd22: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_vscan0_w;
			end
			5'd23: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_base3_w;
			end
			5'd24: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_base2_w;
			end
			5'd25: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_base1_w;
			end
			5'd26: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_base0_w;
			end
			5'd27: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_length3_w;
			end
			5'd28: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_length2_w;
			end
			5'd29: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_length1_w;
			end
			5'd30: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_initiator_length0_w;
			end
			5'd31: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_dma_delay_base3_w;
			end
			6'd32: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_dma_delay_base2_w;
			end
			6'd33: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_dma_delay_base1_w;
			end
			6'd34: begin
				vns_videooverlaysoc_interface3_bank_bus_dat_r <= vns_videooverlaysoc_csrbank3_dma_delay_base0_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank3_underflow_enable0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_underflow_enable_storage_full <= vns_videooverlaysoc_csrbank3_underflow_enable0_r;
	end
	soc_videooverlaysoc_hdmi_core_out0_underflow_enable_re <= vns_videooverlaysoc_csrbank3_underflow_enable0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_enable0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_enable_storage_full <= vns_videooverlaysoc_csrbank3_initiator_enable0_r;
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_enable_re <= vns_videooverlaysoc_csrbank3_initiator_enable0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_hres1_re) begin
		vns_videooverlaysoc_csrbank3_initiator_hres_backstore[3:0] <= vns_videooverlaysoc_csrbank3_initiator_hres1_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_hres0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_storage_full <= {vns_videooverlaysoc_csrbank3_initiator_hres_backstore, vns_videooverlaysoc_csrbank3_initiator_hres0_r};
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_re <= vns_videooverlaysoc_csrbank3_initiator_hres0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_hsync_start1_re) begin
		vns_videooverlaysoc_csrbank3_initiator_hsync_start_backstore[3:0] <= vns_videooverlaysoc_csrbank3_initiator_hsync_start1_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_hsync_start0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_storage_full <= {vns_videooverlaysoc_csrbank3_initiator_hsync_start_backstore, vns_videooverlaysoc_csrbank3_initiator_hsync_start0_r};
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_re <= vns_videooverlaysoc_csrbank3_initiator_hsync_start0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_hsync_end1_re) begin
		vns_videooverlaysoc_csrbank3_initiator_hsync_end_backstore[3:0] <= vns_videooverlaysoc_csrbank3_initiator_hsync_end1_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_hsync_end0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_storage_full <= {vns_videooverlaysoc_csrbank3_initiator_hsync_end_backstore, vns_videooverlaysoc_csrbank3_initiator_hsync_end0_r};
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_re <= vns_videooverlaysoc_csrbank3_initiator_hsync_end0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_hscan1_re) begin
		vns_videooverlaysoc_csrbank3_initiator_hscan_backstore[3:0] <= vns_videooverlaysoc_csrbank3_initiator_hscan1_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_hscan0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_storage_full <= {vns_videooverlaysoc_csrbank3_initiator_hscan_backstore, vns_videooverlaysoc_csrbank3_initiator_hscan0_r};
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_re <= vns_videooverlaysoc_csrbank3_initiator_hscan0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_vres1_re) begin
		vns_videooverlaysoc_csrbank3_initiator_vres_backstore[3:0] <= vns_videooverlaysoc_csrbank3_initiator_vres1_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_vres0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_storage_full <= {vns_videooverlaysoc_csrbank3_initiator_vres_backstore, vns_videooverlaysoc_csrbank3_initiator_vres0_r};
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_re <= vns_videooverlaysoc_csrbank3_initiator_vres0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_vsync_start1_re) begin
		vns_videooverlaysoc_csrbank3_initiator_vsync_start_backstore[3:0] <= vns_videooverlaysoc_csrbank3_initiator_vsync_start1_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_vsync_start0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_storage_full <= {vns_videooverlaysoc_csrbank3_initiator_vsync_start_backstore, vns_videooverlaysoc_csrbank3_initiator_vsync_start0_r};
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_re <= vns_videooverlaysoc_csrbank3_initiator_vsync_start0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_vsync_end1_re) begin
		vns_videooverlaysoc_csrbank3_initiator_vsync_end_backstore[3:0] <= vns_videooverlaysoc_csrbank3_initiator_vsync_end1_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_vsync_end0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_storage_full <= {vns_videooverlaysoc_csrbank3_initiator_vsync_end_backstore, vns_videooverlaysoc_csrbank3_initiator_vsync_end0_r};
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_re <= vns_videooverlaysoc_csrbank3_initiator_vsync_end0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_vscan1_re) begin
		vns_videooverlaysoc_csrbank3_initiator_vscan_backstore[3:0] <= vns_videooverlaysoc_csrbank3_initiator_vscan1_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_vscan0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_storage_full <= {vns_videooverlaysoc_csrbank3_initiator_vscan_backstore, vns_videooverlaysoc_csrbank3_initiator_vscan0_r};
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_re <= vns_videooverlaysoc_csrbank3_initiator_vscan0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_base3_re) begin
		vns_videooverlaysoc_csrbank3_initiator_base_backstore[23:16] <= vns_videooverlaysoc_csrbank3_initiator_base3_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_base2_re) begin
		vns_videooverlaysoc_csrbank3_initiator_base_backstore[15:8] <= vns_videooverlaysoc_csrbank3_initiator_base2_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_base1_re) begin
		vns_videooverlaysoc_csrbank3_initiator_base_backstore[7:0] <= vns_videooverlaysoc_csrbank3_initiator_base1_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_base0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage_full <= {vns_videooverlaysoc_csrbank3_initiator_base_backstore, vns_videooverlaysoc_csrbank3_initiator_base0_r};
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_re <= vns_videooverlaysoc_csrbank3_initiator_base0_re;
	if (vns_videooverlaysoc_csrbank3_initiator_length3_re) begin
		vns_videooverlaysoc_csrbank3_initiator_length_backstore[23:16] <= vns_videooverlaysoc_csrbank3_initiator_length3_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_length2_re) begin
		vns_videooverlaysoc_csrbank3_initiator_length_backstore[15:8] <= vns_videooverlaysoc_csrbank3_initiator_length2_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_length1_re) begin
		vns_videooverlaysoc_csrbank3_initiator_length_backstore[7:0] <= vns_videooverlaysoc_csrbank3_initiator_length1_r;
	end
	if (vns_videooverlaysoc_csrbank3_initiator_length0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage_full <= {vns_videooverlaysoc_csrbank3_initiator_length_backstore, vns_videooverlaysoc_csrbank3_initiator_length0_r};
	end
	soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_re <= vns_videooverlaysoc_csrbank3_initiator_length0_re;
	if (vns_videooverlaysoc_csrbank3_dma_delay_base3_re) begin
		soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full[31:24] <= vns_videooverlaysoc_csrbank3_dma_delay_base3_r;
	end
	if (vns_videooverlaysoc_csrbank3_dma_delay_base2_re) begin
		soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full[23:16] <= vns_videooverlaysoc_csrbank3_dma_delay_base2_r;
	end
	if (vns_videooverlaysoc_csrbank3_dma_delay_base1_re) begin
		soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full[15:8] <= vns_videooverlaysoc_csrbank3_dma_delay_base1_r;
	end
	if (vns_videooverlaysoc_csrbank3_dma_delay_base0_re) begin
		soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full[7:0] <= vns_videooverlaysoc_csrbank3_dma_delay_base0_r;
	end
	soc_videooverlaysoc_hdmi_core_out0_dmareader_re <= vns_videooverlaysoc_csrbank3_dma_delay_base0_re;
	vns_videooverlaysoc_sram0_sel_r <= vns_videooverlaysoc_sram0_sel;
	vns_videooverlaysoc_interface4_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank4_sel) begin
		case (vns_videooverlaysoc_interface4_bank_bus_adr[5:0])
			1'd0: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_edid_hpd_notif_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_edid_hpd_en0_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_mmcm_reset0_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_locked_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_mmcm_read_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_mmcm_write_w;
			end
			3'd6: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_w;
			end
			3'd7: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_mmcm_adr0_w;
			end
			4'd8: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w1_w;
			end
			4'd9: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w0_w;
			end
			4'd10: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r1_w;
			end
			4'd11: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_r0_w;
			end
			4'd12: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_mmcm_write_o_w;
			end
			4'd13: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_mmcm_read_o_w;
			end
			4'd14: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r1_w;
			end
			4'd15: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_o_r0_w;
			end
			5'd16: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_clocking_mmcm_drdy_o_w;
			end
			5'd17: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_dly_ctl_w;
			end
			5'd18: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data0_cap_phase_w;
			end
			5'd19: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture0_phase_reset_w;
			end
			5'd20: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data0_charsync_char_synced_w;
			end
			5'd21: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data0_charsync_ctl_pos_w;
			end
			5'd22: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_wer0_update_w;
			end
			5'd23: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data0_wer_value2_w;
			end
			5'd24: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data0_wer_value1_w;
			end
			5'd25: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data0_wer_value0_w;
			end
			5'd26: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_dly_ctl_w;
			end
			5'd27: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data1_cap_phase_w;
			end
			5'd28: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture1_phase_reset_w;
			end
			5'd29: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data1_charsync_char_synced_w;
			end
			5'd30: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data1_charsync_ctl_pos_w;
			end
			5'd31: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_wer1_update_w;
			end
			6'd32: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data1_wer_value2_w;
			end
			6'd33: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data1_wer_value1_w;
			end
			6'd34: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data1_wer_value0_w;
			end
			6'd35: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_dly_ctl_w;
			end
			6'd36: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data2_cap_phase_w;
			end
			6'd37: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_s7datacapture2_phase_reset_w;
			end
			6'd38: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data2_charsync_char_synced_w;
			end
			6'd39: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data2_charsync_ctl_pos_w;
			end
			6'd40: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in0_wer2_update_w;
			end
			6'd41: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data2_wer_value2_w;
			end
			6'd42: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data2_wer_value1_w;
			end
			6'd43: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_data2_wer_value0_w;
			end
			6'd44: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_chansync_channels_synced_w;
			end
			6'd45: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_decode_terc4_dvimode0_w;
			end
			6'd46: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_resdetection_hres1_w;
			end
			6'd47: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_resdetection_hres0_w;
			end
			6'd48: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_resdetection_vres1_w;
			end
			6'd49: begin
				vns_videooverlaysoc_interface4_bank_bus_dat_r <= vns_videooverlaysoc_csrbank4_resdetection_vres0_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank4_edid_hpd_en0_re) begin
		soc_videooverlaysoc_hdmi_in0_edid_storage_full <= vns_videooverlaysoc_csrbank4_edid_hpd_en0_r;
	end
	soc_videooverlaysoc_hdmi_in0_edid_re <= vns_videooverlaysoc_csrbank4_edid_hpd_en0_re;
	if (vns_videooverlaysoc_csrbank4_clocking_mmcm_reset0_re) begin
		soc_videooverlaysoc_hdmi_in0_mmcm_reset_storage_full <= vns_videooverlaysoc_csrbank4_clocking_mmcm_reset0_r;
	end
	soc_videooverlaysoc_hdmi_in0_mmcm_reset_re <= vns_videooverlaysoc_csrbank4_clocking_mmcm_reset0_re;
	if (vns_videooverlaysoc_csrbank4_clocking_mmcm_adr0_re) begin
		soc_videooverlaysoc_hdmi_in0_mmcm_adr_storage_full[6:0] <= vns_videooverlaysoc_csrbank4_clocking_mmcm_adr0_r;
	end
	soc_videooverlaysoc_hdmi_in0_mmcm_adr_re <= vns_videooverlaysoc_csrbank4_clocking_mmcm_adr0_re;
	if (vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w1_re) begin
		soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage_full[15:8] <= vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w1_r;
	end
	if (vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w0_re) begin
		soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage_full[7:0] <= vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w0_r;
	end
	soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_re <= vns_videooverlaysoc_csrbank4_clocking_mmcm_dat_w0_re;
	if (vns_videooverlaysoc_csrbank4_decode_terc4_dvimode0_re) begin
		soc_videooverlaysoc_hdmi_in0_decode_terc4_storage_full <= vns_videooverlaysoc_csrbank4_decode_terc4_dvimode0_r;
	end
	soc_videooverlaysoc_hdmi_in0_decode_terc4_re <= vns_videooverlaysoc_csrbank4_decode_terc4_dvimode0_re;
	vns_videooverlaysoc_interface5_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank5_sel) begin
		case (vns_videooverlaysoc_interface5_bank_bus_adr[1:0])
			1'd0: begin
				vns_videooverlaysoc_interface5_bank_bus_dat_r <= vns_videooverlaysoc_csrbank5_value3_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface5_bank_bus_dat_r <= vns_videooverlaysoc_csrbank5_value2_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface5_bank_bus_dat_r <= vns_videooverlaysoc_csrbank5_value1_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface5_bank_bus_dat_r <= vns_videooverlaysoc_csrbank5_value0_w;
			end
		endcase
	end
	vns_videooverlaysoc_sram1_sel_r <= vns_videooverlaysoc_sram1_sel;
	vns_videooverlaysoc_interface6_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank6_sel) begin
		case (vns_videooverlaysoc_interface6_bank_bus_adr[5:0])
			1'd0: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_edid_hpd_notif_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_edid_hpd_en0_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_clocking_mmcm_reset0_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_clocking_locked_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_mmcm_read_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_mmcm_write_w;
			end
			3'd6: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_clocking_mmcm_drdy_w;
			end
			3'd7: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_clocking_mmcm_adr0_w;
			end
			4'd8: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w1_w;
			end
			4'd9: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w0_w;
			end
			4'd10: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r1_w;
			end
			4'd11: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_r0_w;
			end
			4'd12: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_dly_ctl_w;
			end
			4'd13: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data0_cap_phase_w;
			end
			4'd14: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture0_phase_reset_w;
			end
			4'd15: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data0_charsync_char_synced_w;
			end
			5'd16: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data0_charsync_ctl_pos_w;
			end
			5'd17: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_wer0_update_w;
			end
			5'd18: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data0_wer_value2_w;
			end
			5'd19: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data0_wer_value1_w;
			end
			5'd20: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data0_wer_value0_w;
			end
			5'd21: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_dly_ctl_w;
			end
			5'd22: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data1_cap_phase_w;
			end
			5'd23: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture1_phase_reset_w;
			end
			5'd24: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data1_charsync_char_synced_w;
			end
			5'd25: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data1_charsync_ctl_pos_w;
			end
			5'd26: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_wer1_update_w;
			end
			5'd27: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data1_wer_value2_w;
			end
			5'd28: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data1_wer_value1_w;
			end
			5'd29: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data1_wer_value0_w;
			end
			5'd30: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_dly_ctl_w;
			end
			5'd31: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data2_cap_phase_w;
			end
			6'd32: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_s7datacapture2_phase_reset_w;
			end
			6'd33: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data2_charsync_char_synced_w;
			end
			6'd34: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data2_charsync_ctl_pos_w;
			end
			6'd35: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_wer2_update_w;
			end
			6'd36: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data2_wer_value2_w;
			end
			6'd37: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data2_wer_value1_w;
			end
			6'd38: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_data2_wer_value0_w;
			end
			6'd39: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_chansync_channels_synced_w;
			end
			6'd40: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_decode_terc4_dvimode0_w;
			end
			6'd41: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_resdetection_hres1_w;
			end
			6'd42: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_resdetection_hres0_w;
			end
			6'd43: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_resdetection_vres1_w;
			end
			6'd44: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_resdetection_vres0_w;
			end
			6'd45: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_frame_overflow_w;
			end
			6'd46: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_frame_size3_w;
			end
			6'd47: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_frame_size2_w;
			end
			6'd48: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_frame_size1_w;
			end
			6'd49: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_frame_size0_w;
			end
			6'd50: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_slot0_status0_w;
			end
			6'd51: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_slot0_address3_w;
			end
			6'd52: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_slot0_address2_w;
			end
			6'd53: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_slot0_address1_w;
			end
			6'd54: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_slot0_address0_w;
			end
			6'd55: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_slot1_status0_w;
			end
			6'd56: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_slot1_address3_w;
			end
			6'd57: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_slot1_address2_w;
			end
			6'd58: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_slot1_address1_w;
			end
			6'd59: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_slot1_address0_w;
			end
			6'd60: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_status_w;
			end
			6'd61: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= soc_videooverlaysoc_hdmi_in1_dma_slot_array_pending_w;
			end
			6'd62: begin
				vns_videooverlaysoc_interface6_bank_bus_dat_r <= vns_videooverlaysoc_csrbank6_dma_ev_enable0_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank6_edid_hpd_en0_re) begin
		soc_videooverlaysoc_hdmi_in1_edid_storage_full <= vns_videooverlaysoc_csrbank6_edid_hpd_en0_r;
	end
	soc_videooverlaysoc_hdmi_in1_edid_re <= vns_videooverlaysoc_csrbank6_edid_hpd_en0_re;
	if (vns_videooverlaysoc_csrbank6_clocking_mmcm_reset0_re) begin
		soc_videooverlaysoc_hdmi_in1_mmcm_reset_storage_full <= vns_videooverlaysoc_csrbank6_clocking_mmcm_reset0_r;
	end
	soc_videooverlaysoc_hdmi_in1_mmcm_reset_re <= vns_videooverlaysoc_csrbank6_clocking_mmcm_reset0_re;
	if (vns_videooverlaysoc_csrbank6_clocking_mmcm_adr0_re) begin
		soc_videooverlaysoc_hdmi_in1_mmcm_adr_storage_full[6:0] <= vns_videooverlaysoc_csrbank6_clocking_mmcm_adr0_r;
	end
	soc_videooverlaysoc_hdmi_in1_mmcm_adr_re <= vns_videooverlaysoc_csrbank6_clocking_mmcm_adr0_re;
	if (vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w1_re) begin
		soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_storage_full[15:8] <= vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w1_r;
	end
	if (vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w0_re) begin
		soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_storage_full[7:0] <= vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w0_r;
	end
	soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_re <= vns_videooverlaysoc_csrbank6_clocking_mmcm_dat_w0_re;
	if (vns_videooverlaysoc_csrbank6_decode_terc4_dvimode0_re) begin
		soc_videooverlaysoc_hdmi_in1_decode_terc4_storage_full <= vns_videooverlaysoc_csrbank6_decode_terc4_dvimode0_r;
	end
	soc_videooverlaysoc_hdmi_in1_decode_terc4_re <= vns_videooverlaysoc_csrbank6_decode_terc4_dvimode0_re;
	if (vns_videooverlaysoc_csrbank6_dma_frame_size3_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full[28:24] <= vns_videooverlaysoc_csrbank6_dma_frame_size3_r;
	end
	if (vns_videooverlaysoc_csrbank6_dma_frame_size2_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full[23:16] <= vns_videooverlaysoc_csrbank6_dma_frame_size2_r;
	end
	if (vns_videooverlaysoc_csrbank6_dma_frame_size1_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full[15:8] <= vns_videooverlaysoc_csrbank6_dma_frame_size1_r;
	end
	if (vns_videooverlaysoc_csrbank6_dma_frame_size0_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full[7:0] <= vns_videooverlaysoc_csrbank6_dma_frame_size0_r;
	end
	soc_videooverlaysoc_hdmi_in1_dma_frame_size_re <= vns_videooverlaysoc_csrbank6_dma_frame_size0_re;
	if (soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_we) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_storage_full <= (soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_dat_w <<< 1'd0);
	end
	if (vns_videooverlaysoc_csrbank6_dma_slot0_status0_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_storage_full[1:0] <= vns_videooverlaysoc_csrbank6_dma_slot0_status0_r;
	end
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_re <= vns_videooverlaysoc_csrbank6_dma_slot0_status0_re;
	if (soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_we) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full <= (soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_dat_w <<< 3'd5);
	end
	if (vns_videooverlaysoc_csrbank6_dma_slot0_address3_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[28:24] <= vns_videooverlaysoc_csrbank6_dma_slot0_address3_r;
	end
	if (vns_videooverlaysoc_csrbank6_dma_slot0_address2_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[23:16] <= vns_videooverlaysoc_csrbank6_dma_slot0_address2_r;
	end
	if (vns_videooverlaysoc_csrbank6_dma_slot0_address1_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[15:8] <= vns_videooverlaysoc_csrbank6_dma_slot0_address1_r;
	end
	if (vns_videooverlaysoc_csrbank6_dma_slot0_address0_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[7:0] <= vns_videooverlaysoc_csrbank6_dma_slot0_address0_r;
	end
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_re <= vns_videooverlaysoc_csrbank6_dma_slot0_address0_re;
	if (soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_we) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_storage_full <= (soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_dat_w <<< 1'd0);
	end
	if (vns_videooverlaysoc_csrbank6_dma_slot1_status0_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_storage_full[1:0] <= vns_videooverlaysoc_csrbank6_dma_slot1_status0_r;
	end
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_re <= vns_videooverlaysoc_csrbank6_dma_slot1_status0_re;
	if (soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_we) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full <= (soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_dat_w <<< 3'd5);
	end
	if (vns_videooverlaysoc_csrbank6_dma_slot1_address3_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[28:24] <= vns_videooverlaysoc_csrbank6_dma_slot1_address3_r;
	end
	if (vns_videooverlaysoc_csrbank6_dma_slot1_address2_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[23:16] <= vns_videooverlaysoc_csrbank6_dma_slot1_address2_r;
	end
	if (vns_videooverlaysoc_csrbank6_dma_slot1_address1_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[15:8] <= vns_videooverlaysoc_csrbank6_dma_slot1_address1_r;
	end
	if (vns_videooverlaysoc_csrbank6_dma_slot1_address0_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[7:0] <= vns_videooverlaysoc_csrbank6_dma_slot1_address0_r;
	end
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_re <= vns_videooverlaysoc_csrbank6_dma_slot1_address0_re;
	if (vns_videooverlaysoc_csrbank6_dma_ev_enable0_re) begin
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_storage_full[1:0] <= vns_videooverlaysoc_csrbank6_dma_ev_enable0_r;
	end
	soc_videooverlaysoc_hdmi_in1_dma_slot_array_re <= vns_videooverlaysoc_csrbank6_dma_ev_enable0_re;
	vns_videooverlaysoc_interface7_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank7_sel) begin
		case (vns_videooverlaysoc_interface7_bank_bus_adr[1:0])
			1'd0: begin
				vns_videooverlaysoc_interface7_bank_bus_dat_r <= vns_videooverlaysoc_csrbank7_value3_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface7_bank_bus_dat_r <= vns_videooverlaysoc_csrbank7_value2_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface7_bank_bus_dat_r <= vns_videooverlaysoc_csrbank7_value1_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface7_bank_bus_dat_r <= vns_videooverlaysoc_csrbank7_value0_w;
			end
		endcase
	end
	vns_videooverlaysoc_interface8_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank8_sel) begin
		case (vns_videooverlaysoc_interface8_bank_bus_adr[0])
			1'd0: begin
				vns_videooverlaysoc_interface8_bank_bus_dat_r <= vns_videooverlaysoc_csrbank8_edid_snoop_adr0_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface8_bank_bus_dat_r <= vns_videooverlaysoc_csrbank8_edid_snoop_dat_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank8_edid_snoop_adr0_re) begin
		soc_videooverlaysoc_i2c_snoop_storage_full[7:0] <= vns_videooverlaysoc_csrbank8_edid_snoop_adr0_r;
	end
	soc_videooverlaysoc_i2c_snoop_re <= vns_videooverlaysoc_csrbank8_edid_snoop_adr0_re;
	vns_videooverlaysoc_sram2_sel_r <= vns_videooverlaysoc_sram2_sel;
	vns_videooverlaysoc_interface9_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank9_sel) begin
		case (vns_videooverlaysoc_interface9_bank_bus_adr[3:0])
			1'd0: begin
				vns_videooverlaysoc_interface9_bank_bus_dat_r <= vns_videooverlaysoc_csrbank9_hrect_start1_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface9_bank_bus_dat_r <= vns_videooverlaysoc_csrbank9_hrect_start0_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface9_bank_bus_dat_r <= vns_videooverlaysoc_csrbank9_hrect_end1_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface9_bank_bus_dat_r <= vns_videooverlaysoc_csrbank9_hrect_end0_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface9_bank_bus_dat_r <= vns_videooverlaysoc_csrbank9_vrect_start1_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface9_bank_bus_dat_r <= vns_videooverlaysoc_csrbank9_vrect_start0_w;
			end
			3'd6: begin
				vns_videooverlaysoc_interface9_bank_bus_dat_r <= vns_videooverlaysoc_csrbank9_vrect_end1_w;
			end
			3'd7: begin
				vns_videooverlaysoc_interface9_bank_bus_dat_r <= vns_videooverlaysoc_csrbank9_vrect_end0_w;
			end
			4'd8: begin
				vns_videooverlaysoc_interface9_bank_bus_dat_r <= vns_videooverlaysoc_csrbank9_rect_thresh0_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank9_hrect_start1_re) begin
		soc_videooverlaysoc_hrect_start_storage_full[11:8] <= vns_videooverlaysoc_csrbank9_hrect_start1_r;
	end
	if (vns_videooverlaysoc_csrbank9_hrect_start0_re) begin
		soc_videooverlaysoc_hrect_start_storage_full[7:0] <= vns_videooverlaysoc_csrbank9_hrect_start0_r;
	end
	soc_videooverlaysoc_hrect_start_re <= vns_videooverlaysoc_csrbank9_hrect_start0_re;
	if (vns_videooverlaysoc_csrbank9_hrect_end1_re) begin
		soc_videooverlaysoc_hrect_end_storage_full[11:8] <= vns_videooverlaysoc_csrbank9_hrect_end1_r;
	end
	if (vns_videooverlaysoc_csrbank9_hrect_end0_re) begin
		soc_videooverlaysoc_hrect_end_storage_full[7:0] <= vns_videooverlaysoc_csrbank9_hrect_end0_r;
	end
	soc_videooverlaysoc_hrect_end_re <= vns_videooverlaysoc_csrbank9_hrect_end0_re;
	if (vns_videooverlaysoc_csrbank9_vrect_start1_re) begin
		soc_videooverlaysoc_vrect_start_storage_full[11:8] <= vns_videooverlaysoc_csrbank9_vrect_start1_r;
	end
	if (vns_videooverlaysoc_csrbank9_vrect_start0_re) begin
		soc_videooverlaysoc_vrect_start_storage_full[7:0] <= vns_videooverlaysoc_csrbank9_vrect_start0_r;
	end
	soc_videooverlaysoc_vrect_start_re <= vns_videooverlaysoc_csrbank9_vrect_start0_re;
	if (vns_videooverlaysoc_csrbank9_vrect_end1_re) begin
		soc_videooverlaysoc_vrect_end_storage_full[11:8] <= vns_videooverlaysoc_csrbank9_vrect_end1_r;
	end
	if (vns_videooverlaysoc_csrbank9_vrect_end0_re) begin
		soc_videooverlaysoc_vrect_end_storage_full[7:0] <= vns_videooverlaysoc_csrbank9_vrect_end0_r;
	end
	soc_videooverlaysoc_vrect_end_re <= vns_videooverlaysoc_csrbank9_vrect_end0_re;
	if (vns_videooverlaysoc_csrbank9_rect_thresh0_re) begin
		soc_videooverlaysoc_rect_thresh_storage_full[7:0] <= vns_videooverlaysoc_csrbank9_rect_thresh0_r;
	end
	soc_videooverlaysoc_rect_thresh_re <= vns_videooverlaysoc_csrbank9_rect_thresh0_re;
	vns_videooverlaysoc_interface10_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank10_sel) begin
		case (vns_videooverlaysoc_interface10_bank_bus_adr[6:0])
			1'd0: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_control0_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_command0_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_issue_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_address1_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_address0_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_baddress0_w;
			end
			3'd6: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata7_w;
			end
			3'd7: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata6_w;
			end
			4'd8: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata5_w;
			end
			4'd9: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata4_w;
			end
			4'd10: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata3_w;
			end
			4'd11: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata2_w;
			end
			4'd12: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata1_w;
			end
			4'd13: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata0_w;
			end
			4'd14: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_rddata7_w;
			end
			4'd15: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_rddata6_w;
			end
			5'd16: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_rddata5_w;
			end
			5'd17: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_rddata4_w;
			end
			5'd18: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_rddata3_w;
			end
			5'd19: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_rddata2_w;
			end
			5'd20: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_rddata1_w;
			end
			5'd21: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi0_rddata0_w;
			end
			5'd22: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_command0_w;
			end
			5'd23: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_issue_w;
			end
			5'd24: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_address1_w;
			end
			5'd25: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_address0_w;
			end
			5'd26: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_baddress0_w;
			end
			5'd27: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata7_w;
			end
			5'd28: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata6_w;
			end
			5'd29: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata5_w;
			end
			5'd30: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata4_w;
			end
			5'd31: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata3_w;
			end
			6'd32: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata2_w;
			end
			6'd33: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata1_w;
			end
			6'd34: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata0_w;
			end
			6'd35: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_rddata7_w;
			end
			6'd36: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_rddata6_w;
			end
			6'd37: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_rddata5_w;
			end
			6'd38: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_rddata4_w;
			end
			6'd39: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_rddata3_w;
			end
			6'd40: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_rddata2_w;
			end
			6'd41: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_rddata1_w;
			end
			6'd42: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi1_rddata0_w;
			end
			6'd43: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_command0_w;
			end
			6'd44: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_issue_w;
			end
			6'd45: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_address1_w;
			end
			6'd46: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_address0_w;
			end
			6'd47: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_baddress0_w;
			end
			6'd48: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata7_w;
			end
			6'd49: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata6_w;
			end
			6'd50: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata5_w;
			end
			6'd51: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata4_w;
			end
			6'd52: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata3_w;
			end
			6'd53: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata2_w;
			end
			6'd54: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata1_w;
			end
			6'd55: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata0_w;
			end
			6'd56: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_rddata7_w;
			end
			6'd57: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_rddata6_w;
			end
			6'd58: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_rddata5_w;
			end
			6'd59: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_rddata4_w;
			end
			6'd60: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_rddata3_w;
			end
			6'd61: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_rddata2_w;
			end
			6'd62: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_rddata1_w;
			end
			6'd63: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi2_rddata0_w;
			end
			7'd64: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_command0_w;
			end
			7'd65: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_issue_w;
			end
			7'd66: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_address1_w;
			end
			7'd67: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_address0_w;
			end
			7'd68: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_baddress0_w;
			end
			7'd69: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata7_w;
			end
			7'd70: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata6_w;
			end
			7'd71: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata5_w;
			end
			7'd72: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata4_w;
			end
			7'd73: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata3_w;
			end
			7'd74: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata2_w;
			end
			7'd75: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata1_w;
			end
			7'd76: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata0_w;
			end
			7'd77: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_rddata7_w;
			end
			7'd78: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_rddata6_w;
			end
			7'd79: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_rddata5_w;
			end
			7'd80: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_rddata4_w;
			end
			7'd81: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_rddata3_w;
			end
			7'd82: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_rddata2_w;
			end
			7'd83: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_rddata1_w;
			end
			7'd84: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_dfii_pi3_rddata0_w;
			end
			7'd85: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_update_w;
			end
			7'd86: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads2_w;
			end
			7'd87: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads1_w;
			end
			7'd88: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_controller_bandwidth_nreads0_w;
			end
			7'd89: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites2_w;
			end
			7'd90: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites1_w;
			end
			7'd91: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_controller_bandwidth_nwrites0_w;
			end
			7'd92: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width1_w;
			end
			7'd93: begin
				vns_videooverlaysoc_interface10_bank_bus_dat_r <= vns_videooverlaysoc_csrbank10_controller_bandwidth_data_width0_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank10_dfii_control0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_storage_full[3:0] <= vns_videooverlaysoc_csrbank10_dfii_control0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_re <= vns_videooverlaysoc_csrbank10_dfii_control0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_command0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage_full[5:0] <= vns_videooverlaysoc_csrbank10_dfii_pi0_command0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_re <= vns_videooverlaysoc_csrbank10_dfii_pi0_command0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_address1_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_storage_full[13:8] <= vns_videooverlaysoc_csrbank10_dfii_pi0_address1_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_address0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_storage_full[7:0] <= vns_videooverlaysoc_csrbank10_dfii_pi0_address0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_re <= vns_videooverlaysoc_csrbank10_dfii_pi0_address0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_baddress0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_storage_full[2:0] <= vns_videooverlaysoc_csrbank10_dfii_pi0_baddress0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_re <= vns_videooverlaysoc_csrbank10_dfii_pi0_baddress0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata7_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[63:56] <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata7_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata6_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[55:48] <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata6_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata5_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[47:40] <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata5_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata4_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[39:32] <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata4_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata3_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[31:24] <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata3_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata2_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[23:16] <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata2_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata1_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[15:8] <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata1_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full[7:0] <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_re <= vns_videooverlaysoc_csrbank10_dfii_pi0_wrdata0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_command0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage_full[5:0] <= vns_videooverlaysoc_csrbank10_dfii_pi1_command0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_re <= vns_videooverlaysoc_csrbank10_dfii_pi1_command0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_address1_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_storage_full[13:8] <= vns_videooverlaysoc_csrbank10_dfii_pi1_address1_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_address0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_storage_full[7:0] <= vns_videooverlaysoc_csrbank10_dfii_pi1_address0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_re <= vns_videooverlaysoc_csrbank10_dfii_pi1_address0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_baddress0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_storage_full[2:0] <= vns_videooverlaysoc_csrbank10_dfii_pi1_baddress0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_re <= vns_videooverlaysoc_csrbank10_dfii_pi1_baddress0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata7_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[63:56] <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata7_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata6_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[55:48] <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata6_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata5_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[47:40] <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata5_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata4_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[39:32] <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata4_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata3_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[31:24] <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata3_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata2_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[23:16] <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata2_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata1_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[15:8] <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata1_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full[7:0] <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_re <= vns_videooverlaysoc_csrbank10_dfii_pi1_wrdata0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_command0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage_full[5:0] <= vns_videooverlaysoc_csrbank10_dfii_pi2_command0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_re <= vns_videooverlaysoc_csrbank10_dfii_pi2_command0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_address1_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_storage_full[13:8] <= vns_videooverlaysoc_csrbank10_dfii_pi2_address1_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_address0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_storage_full[7:0] <= vns_videooverlaysoc_csrbank10_dfii_pi2_address0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_re <= vns_videooverlaysoc_csrbank10_dfii_pi2_address0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_baddress0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_storage_full[2:0] <= vns_videooverlaysoc_csrbank10_dfii_pi2_baddress0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_re <= vns_videooverlaysoc_csrbank10_dfii_pi2_baddress0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata7_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[63:56] <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata7_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata6_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[55:48] <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata6_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata5_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[47:40] <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata5_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata4_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[39:32] <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata4_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata3_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[31:24] <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata3_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata2_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[23:16] <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata2_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata1_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[15:8] <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata1_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full[7:0] <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_re <= vns_videooverlaysoc_csrbank10_dfii_pi2_wrdata0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_command0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage_full[5:0] <= vns_videooverlaysoc_csrbank10_dfii_pi3_command0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_re <= vns_videooverlaysoc_csrbank10_dfii_pi3_command0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_address1_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_storage_full[13:8] <= vns_videooverlaysoc_csrbank10_dfii_pi3_address1_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_address0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_storage_full[7:0] <= vns_videooverlaysoc_csrbank10_dfii_pi3_address0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_re <= vns_videooverlaysoc_csrbank10_dfii_pi3_address0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_baddress0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_storage_full[2:0] <= vns_videooverlaysoc_csrbank10_dfii_pi3_baddress0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_re <= vns_videooverlaysoc_csrbank10_dfii_pi3_baddress0_re;
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata7_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[63:56] <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata7_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata6_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[55:48] <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata6_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata5_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[47:40] <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata5_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata4_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[39:32] <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata4_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata3_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[31:24] <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata3_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata2_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[23:16] <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata2_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata1_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[15:8] <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata1_r;
	end
	if (vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata0_re) begin
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full[7:0] <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_re <= vns_videooverlaysoc_csrbank10_dfii_pi3_wrdata0_re;
	vns_videooverlaysoc_interface11_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank11_sel) begin
		case (vns_videooverlaysoc_interface11_bank_bus_adr[4:0])
			1'd0: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_load3_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_load2_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_load1_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_load0_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_reload3_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_reload2_w;
			end
			3'd6: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_reload1_w;
			end
			3'd7: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_reload0_w;
			end
			4'd8: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_en0_w;
			end
			4'd9: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_update_value_w;
			end
			4'd10: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_value3_w;
			end
			4'd11: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_value2_w;
			end
			4'd12: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_value1_w;
			end
			4'd13: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_value0_w;
			end
			4'd14: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_status_w;
			end
			4'd15: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_pending_w;
			end
			5'd16: begin
				vns_videooverlaysoc_interface11_bank_bus_dat_r <= vns_videooverlaysoc_csrbank11_ev_enable0_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank11_load3_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full[31:24] <= vns_videooverlaysoc_csrbank11_load3_r;
	end
	if (vns_videooverlaysoc_csrbank11_load2_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full[23:16] <= vns_videooverlaysoc_csrbank11_load2_r;
	end
	if (vns_videooverlaysoc_csrbank11_load1_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full[15:8] <= vns_videooverlaysoc_csrbank11_load1_r;
	end
	if (vns_videooverlaysoc_csrbank11_load0_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full[7:0] <= vns_videooverlaysoc_csrbank11_load0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_re <= vns_videooverlaysoc_csrbank11_load0_re;
	if (vns_videooverlaysoc_csrbank11_reload3_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full[31:24] <= vns_videooverlaysoc_csrbank11_reload3_r;
	end
	if (vns_videooverlaysoc_csrbank11_reload2_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full[23:16] <= vns_videooverlaysoc_csrbank11_reload2_r;
	end
	if (vns_videooverlaysoc_csrbank11_reload1_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full[15:8] <= vns_videooverlaysoc_csrbank11_reload1_r;
	end
	if (vns_videooverlaysoc_csrbank11_reload0_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full[7:0] <= vns_videooverlaysoc_csrbank11_reload0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_re <= vns_videooverlaysoc_csrbank11_reload0_re;
	if (vns_videooverlaysoc_csrbank11_en0_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_storage_full <= vns_videooverlaysoc_csrbank11_en0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_re <= vns_videooverlaysoc_csrbank11_en0_re;
	if (vns_videooverlaysoc_csrbank11_ev_enable0_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_storage_full <= vns_videooverlaysoc_csrbank11_ev_enable0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_re <= vns_videooverlaysoc_csrbank11_ev_enable0_re;
	vns_videooverlaysoc_interface12_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank12_sel) begin
		case (vns_videooverlaysoc_interface12_bank_bus_adr[2:0])
			1'd0: begin
				vns_videooverlaysoc_interface12_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rxtx_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface12_bank_bus_dat_r <= vns_videooverlaysoc_csrbank12_txfull_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface12_bank_bus_dat_r <= vns_videooverlaysoc_csrbank12_rxempty_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface12_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_status_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface12_bank_bus_dat_r <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_pending_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface12_bank_bus_dat_r <= vns_videooverlaysoc_csrbank12_ev_enable0_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank12_ev_enable0_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_storage_full[1:0] <= vns_videooverlaysoc_csrbank12_ev_enable0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_re <= vns_videooverlaysoc_csrbank12_ev_enable0_re;
	vns_videooverlaysoc_interface13_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank13_sel) begin
		case (vns_videooverlaysoc_interface13_bank_bus_adr[1:0])
			1'd0: begin
				vns_videooverlaysoc_interface13_bank_bus_dat_r <= vns_videooverlaysoc_csrbank13_tuning_word3_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface13_bank_bus_dat_r <= vns_videooverlaysoc_csrbank13_tuning_word2_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface13_bank_bus_dat_r <= vns_videooverlaysoc_csrbank13_tuning_word1_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface13_bank_bus_dat_r <= vns_videooverlaysoc_csrbank13_tuning_word0_w;
			end
		endcase
	end
	if (vns_videooverlaysoc_csrbank13_tuning_word3_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full[31:24] <= vns_videooverlaysoc_csrbank13_tuning_word3_r;
	end
	if (vns_videooverlaysoc_csrbank13_tuning_word2_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full[23:16] <= vns_videooverlaysoc_csrbank13_tuning_word2_r;
	end
	if (vns_videooverlaysoc_csrbank13_tuning_word1_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full[15:8] <= vns_videooverlaysoc_csrbank13_tuning_word1_r;
	end
	if (vns_videooverlaysoc_csrbank13_tuning_word0_re) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full[7:0] <= vns_videooverlaysoc_csrbank13_tuning_word0_r;
	end
	soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_re <= vns_videooverlaysoc_csrbank13_tuning_word0_re;
	vns_videooverlaysoc_interface14_bank_bus_dat_r <= 1'd0;
	if (vns_videooverlaysoc_csrbank14_sel) begin
		case (vns_videooverlaysoc_interface14_bank_bus_adr[2:0])
			1'd0: begin
				vns_videooverlaysoc_interface14_bank_bus_dat_r <= vns_videooverlaysoc_csrbank14_temperature1_w;
			end
			1'd1: begin
				vns_videooverlaysoc_interface14_bank_bus_dat_r <= vns_videooverlaysoc_csrbank14_temperature0_w;
			end
			2'd2: begin
				vns_videooverlaysoc_interface14_bank_bus_dat_r <= vns_videooverlaysoc_csrbank14_vccint1_w;
			end
			2'd3: begin
				vns_videooverlaysoc_interface14_bank_bus_dat_r <= vns_videooverlaysoc_csrbank14_vccint0_w;
			end
			3'd4: begin
				vns_videooverlaysoc_interface14_bank_bus_dat_r <= vns_videooverlaysoc_csrbank14_vccaux1_w;
			end
			3'd5: begin
				vns_videooverlaysoc_interface14_bank_bus_dat_r <= vns_videooverlaysoc_csrbank14_vccaux0_w;
			end
			3'd6: begin
				vns_videooverlaysoc_interface14_bank_bus_dat_r <= vns_videooverlaysoc_csrbank14_vccbram1_w;
			end
			3'd7: begin
				vns_videooverlaysoc_interface14_bank_bus_dat_r <= vns_videooverlaysoc_csrbank14_vccbram0_w;
			end
		endcase
	end
	if (sys_rst) begin
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_storage_full <= 32'd305419896;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_ctrl_bus_errors <= 32'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_err <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_d_err <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_cpu_reset <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_valid <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_wr <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_address <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_data <= 32'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_reset_debug_logic <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_complete <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_in_progress <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_transfer_wait_for_ack <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_dat_r <= 32'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_debug_bus_ack <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_bus_ack <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_bus_ack <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_adr <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_we <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_interface_dat_w <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_dat_r <= 32'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_bus_wishbone_ack <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_counter <= 2'd0;
		serial_tx <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_storage_full <= 32'd4947802;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_sink_ready <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_uart_clk_txen <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_phase_accumulator_tx <= 32'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_reg <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_bitcount <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_tx_busy <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_valid <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_source_payload_data <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_uart_clk_rxen <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_phase_accumulator_rx <= 32'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_r <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_reg <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_bitcount <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_phy_rx_busy <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_pending <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_old_trigger <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_pending <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_old_trigger <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_storage_full <= 2'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_eventmanager_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_readable <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_level0 <= 5'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_produce <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_consume <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_readable <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_level0 <= 5'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_produce <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_consume <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_storage_full <= 32'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_load_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_storage_full <= 32'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_reload_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_storage_full <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_en_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value_status <= 32'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_pending <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_zero_old_trigger <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_storage_full <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_eventmanager_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_timer0_value <= 32'd0;
		soc_videooverlaysoc_videooverlaysoc_temperature_status <= 12'd0;
		soc_videooverlaysoc_videooverlaysoc_vccint_status <= 12'd0;
		soc_videooverlaysoc_videooverlaysoc_vccaux_status <= 12'd0;
		soc_videooverlaysoc_videooverlaysoc_vccbram_status <= 12'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_half_sys8x_taps_storage_full <= 4'd8;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_half_sys8x_taps_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage_full <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_rddata_valid <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_rddata_valid <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_rddata_valid <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_rddata_valid <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dqs <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip0_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip1_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip2_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip3_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip4_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip5_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip6_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip7_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip8_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip9_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip10_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip11_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip12_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip13_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip14_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip15_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip16_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip17_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip18_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip19_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip20_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip21_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip22_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip23_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip24_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip25_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip26_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip27_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip28_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip29_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip30_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_o <= 8'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_value <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_bitslip31_r <= 16'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en0 <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en1 <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en2 <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en3 <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en4 <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en5 <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en6 <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_n_rddata_en7 <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_a7ddrphy_last_wrdata_en <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_storage_full <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_storage_full <= 6'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_command_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_storage_full <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_address_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_storage_full <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_baddress_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_storage_full <= 64'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_wrdata_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector0_status <= 64'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_storage_full <= 6'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_command_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_storage_full <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_address_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_storage_full <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_baddress_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_storage_full <= 64'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_wrdata_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector1_status <= 64'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_storage_full <= 6'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_command_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_storage_full <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_address_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_storage_full <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_baddress_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_storage_full <= 64'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_wrdata_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector2_status <= 64'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_storage_full <= 6'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_command_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_storage_full <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_address_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_storage_full <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_baddress_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_storage_full <= 64'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_wrdata_re <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_phaseinjector3_status <= 64'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_address <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_bank <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cas_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_cs_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_ras_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_we_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_wrdata_en <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p0_rddata_en <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_address <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_bank <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cas_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_cs_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_ras_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_we_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_wrdata_en <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p1_rddata_en <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_address <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_bank <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cas_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_cs_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_ras_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_we_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_wrdata_en <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p2_rddata_en <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_address <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_bank <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cas_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_cs_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_ras_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_we_n <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_wrdata_en <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_dfi_p3_rddata_en <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_a <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ba <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_cas <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_ras <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_cmd_payload_we <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_seq_done <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_counter <= 5'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_count <= 10'd782;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_level <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_produce <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_consume <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_we <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_source_payload_addr <= 21'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_valid_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_first_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_last_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_row_opened <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_twtpcon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trccon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_trascon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_level <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_produce <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_consume <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_we <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_source_payload_addr <= 21'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_valid_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_first_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_last_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_row_opened <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_twtpcon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trccon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_trascon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_level <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_produce <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_consume <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_we <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_source_payload_addr <= 21'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_valid_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_first_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_last_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_row_opened <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_twtpcon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trccon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_trascon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_level <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_produce <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_consume <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_we <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_source_payload_addr <= 21'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_valid_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_first_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_last_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_row_opened <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_twtpcon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trccon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_trascon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_level <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_produce <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_consume <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_we <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_source_payload_addr <= 21'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_valid_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_first_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_last_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_row_opened <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_twtpcon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trccon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_trascon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_level <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_produce <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_consume <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_we <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_source_payload_addr <= 21'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_valid_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_first_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_last_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_row_opened <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_twtpcon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trccon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_trascon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_level <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_produce <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_consume <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_we <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_source_payload_addr <= 21'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_valid_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_first_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_last_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_row_opened <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_twtpcon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trccon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_trascon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_level <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_produce <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_consume <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_we <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_source_payload_addr <= 21'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_valid_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_first_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_last_n <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row <= 14'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_row_opened <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_twtpcon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trccon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_trascon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_choose_cmd_grant <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_choose_req_grant <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_trrdcon_count <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_tfawcon_window <= 5'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_tccdcon_count <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_ready <= 1'd1;
		soc_videooverlaysoc_videooverlaysoc_sdram_twtrcon_count <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_time0 <= 5'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_time1 <= 4'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads_status <= 24'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites_status <= 24'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_valid <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_ready <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_is_read <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_cmd_is_write <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_counter <= 24'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_period <= 1'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads <= 24'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites <= 24'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nreads_r <= 24'd0;
		soc_videooverlaysoc_videooverlaysoc_sdram_bandwidth_nwrites_r <= 24'd0;
		soc_videooverlaysoc_videooverlaysoc_adr_offset_r <= 3'd0;
		soc_videooverlaysoc_videooverlaysoc_sys_counter <= 32'd0;
		soc_videooverlaysoc_hdmi_in0_freq_period_counter <= 32'd0;
		soc_videooverlaysoc_hdmi_in0_freq_sampler_o <= 32'd0;
		soc_videooverlaysoc_hdmi_in0_freq_sampler_counter <= 32'd0;
		soc_videooverlaysoc_hdmi_in0_freq_sampler_i_d <= 6'd0;
		soc_videooverlaysoc_hdmi_in0_edid_storage_full <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_edid_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_edid_sda_i <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_edid_sda_drv_reg <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_edid_scl_i <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_edid_samp_count <= 6'd0;
		soc_videooverlaysoc_hdmi_in0_edid_samp_carry <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_edid_scl_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_edid_sda_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_edid_din <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_edid_counter <= 4'd0;
		soc_videooverlaysoc_hdmi_in0_edid_is_read <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_edid_offset_counter <= 8'd0;
		soc_videooverlaysoc_hdmi_in0_edid_data_bit <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_edid_data_drv <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_mmcm_reset_storage_full <= 1'd1;
		soc_videooverlaysoc_hdmi_in0_mmcm_reset_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_mmcm_drdy_status <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_mmcm_adr_storage_full <= 7'd0;
		soc_videooverlaysoc_hdmi_in0_mmcm_adr_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage_full <= 16'd0;
		soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_mmcm_drdy_o_status <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_status <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer0_wer_counter_sys <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_status <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer1_wer_counter_sys <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_status <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_wer2_wer_counter_sys <= 24'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_storage_full <= 1'd0;
		soc_videooverlaysoc_hdmi_in0_decode_terc4_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_freq_period_counter <= 32'd0;
		soc_videooverlaysoc_hdmi_in1_freq_sampler_o <= 32'd0;
		soc_videooverlaysoc_hdmi_in1_freq_sampler_counter <= 32'd0;
		soc_videooverlaysoc_hdmi_in1_freq_sampler_i_d <= 6'd0;
		soc_videooverlaysoc_hdmi_in1_edid_storage_full <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_edid_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_edid_sda_i <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_edid_sda_drv_reg <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_edid_scl_i <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_edid_samp_count <= 6'd0;
		soc_videooverlaysoc_hdmi_in1_edid_samp_carry <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_edid_scl_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_edid_sda_r <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_edid_din <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_edid_counter <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_edid_is_read <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_edid_offset_counter <= 8'd0;
		soc_videooverlaysoc_hdmi_in1_edid_data_bit <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_edid_data_drv <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_mmcm_reset_storage_full <= 1'd1;
		soc_videooverlaysoc_hdmi_in1_mmcm_reset_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_mmcm_drdy_status <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_mmcm_adr_storage_full <= 7'd0;
		soc_videooverlaysoc_hdmi_in1_mmcm_adr_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_storage_full <= 16'd0;
		soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_status <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer0_wer_counter_sys <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_status <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer1_wer_counter_sys <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_status <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_wer2_wer_counter_sys <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_storage_full <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_decode_terc4_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q <= 11'd0;
		soc_videooverlaysoc_hdmi_in1_frame_graycounter1_q_binary <= 11'd0;
		soc_videooverlaysoc_hdmi_in1_frame_overflow_mask <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_dma_frame_size_storage_full <= 29'd0;
		soc_videooverlaysoc_hdmi_in1_dma_frame_size_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_storage_full <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_status_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_storage_full <= 29'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot0_address_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_storage_full <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_status_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_storage_full <= 29'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_slot1_address_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_storage_full <= 2'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_re <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_dma_slot_array_current_slot <= 1'd0;
		soc_videooverlaysoc_hdmi_in1_dma_current_address <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_dma_mwords_remaining <= 24'd0;
		soc_videooverlaysoc_hdmi_in1_dma_fifo_level <= 5'd0;
		soc_videooverlaysoc_hdmi_in1_dma_fifo_produce <= 4'd0;
		soc_videooverlaysoc_hdmi_in1_dma_fifo_consume <= 4'd0;
		soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q <= 3'd0;
		soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter1_q_binary <= 3'd0;
		soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q <= 5'd0;
		soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter0_q_binary <= 5'd0;
		soc_videooverlaysoc_hdmi_core_out0_underflow_enable_storage_full <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_underflow_enable_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q <= 2'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter0_q_binary <= 2'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_enable_storage_full <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_enable_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_storage_full <= 12'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage0_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_storage_full <= 12'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage1_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_storage_full <= 12'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage2_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_storage_full <= 12'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage3_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_storage_full <= 12'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage4_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_storage_full <= 12'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage5_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_storage_full <= 12'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage6_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_storage_full <= 12'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage7_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_storage_full <= 32'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage8_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_storage_full <= 32'd0;
		soc_videooverlaysoc_hdmi_core_out0_initiator_csrstorage9_re <= 1'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_storage_full <= 32'd0;
		soc_videooverlaysoc_hdmi_core_out0_dmareader_re <= 1'd0;
		soc_videooverlaysoc_i2c_snoop_storage_full <= 8'd0;
		soc_videooverlaysoc_i2c_snoop_re <= 1'd0;
		soc_videooverlaysoc_hdcp_Km_storage_full <= 56'd0;
		soc_videooverlaysoc_hdcp_Km_re <= 1'd0;
		soc_videooverlaysoc_hdcp_Km_valid_storage_full <= 1'd0;
		soc_videooverlaysoc_hdcp_Km_valid_re <= 1'd0;
		soc_videooverlaysoc_hdcp_hpd_ena_storage_full <= 1'd0;
		soc_videooverlaysoc_hdcp_hpd_ena_re <= 1'd0;
		soc_videooverlaysoc_hrect_start_storage_full <= 12'd0;
		soc_videooverlaysoc_hrect_start_re <= 1'd0;
		soc_videooverlaysoc_hrect_end_storage_full <= 12'd0;
		soc_videooverlaysoc_hrect_end_re <= 1'd0;
		soc_videooverlaysoc_vrect_start_storage_full <= 12'd0;
		soc_videooverlaysoc_vrect_start_re <= 1'd0;
		soc_videooverlaysoc_vrect_end_storage_full <= 12'd0;
		soc_videooverlaysoc_vrect_end_re <= 1'd0;
		soc_videooverlaysoc_rect_thresh_storage_full <= 8'd0;
		soc_videooverlaysoc_rect_thresh_re <= 1'd0;
		soc_videooverlaysoc_packet_liteethetherbonepacketpacketizer_counter <= 1'd0;
		soc_videooverlaysoc_packet_depacketizer_counter <= 1'd0;
		soc_videooverlaysoc_packet_depacketizer_no_payload <= 1'd0;
		soc_videooverlaysoc_record_depacketizer_counter <= 1'd0;
		soc_videooverlaysoc_record_depacketizer_no_payload <= 1'd0;
		soc_videooverlaysoc_record_receiver_fifo_readable <= 1'd0;
		soc_videooverlaysoc_record_receiver_fifo_level0 <= 3'd0;
		soc_videooverlaysoc_record_receiver_fifo_produce <= 2'd0;
		soc_videooverlaysoc_record_receiver_fifo_consume <= 2'd0;
		soc_videooverlaysoc_record_first <= 1'd1;
		soc_videooverlaysoc_record_sender_source_source_payload_data <= 32'd0;
		soc_videooverlaysoc_record_sender_source_source_param_byte_enable <= 8'd0;
		soc_videooverlaysoc_record_sender_source_source_param_rcount <= 8'd0;
		soc_videooverlaysoc_record_sender_source_source_param_wcount <= 8'd0;
		soc_videooverlaysoc_record_sender_fifo_readable <= 1'd0;
		soc_videooverlaysoc_record_sender_fifo_level0 <= 3'd0;
		soc_videooverlaysoc_record_sender_fifo_produce <= 2'd0;
		soc_videooverlaysoc_record_sender_fifo_consume <= 2'd0;
		soc_videooverlaysoc_record_packetizer_counter <= 1'd0;
		soc_videooverlaysoc_dispatcher_first <= 1'd1;
		soc_videooverlaysoc_dispatcher_ongoing1 <= 1'd0;
		soc_videooverlaysoc_dispatcher_sel_ongoing <= 1'd0;
		soc_videooverlaysoc_grant <= 1'd0;
		soc_videooverlaysoc_status0_first <= 1'd1;
		soc_videooverlaysoc_status0_ongoing1 <= 1'd0;
		soc_videooverlaysoc_status1_first <= 1'd1;
		soc_videooverlaysoc_status1_ongoing1 <= 1'd0;
		soc_videooverlaysoc_wishbone_source_payload_addr <= 32'd0;
		soc_videooverlaysoc_wishbone_source_payload_data <= 32'd0;
		soc_videooverlaysoc_wishbone_source_param_we <= 1'd0;
		soc_videooverlaysoc_wishbone_source_param_count <= 8'd0;
		soc_videooverlaysoc_wishbone_source_param_base_addr <= 32'd0;
		soc_videooverlaysoc_wishbone_source_param_be <= 4'd0;
		fpga_led40 <= 1'd0;
		vns_refresher_state <= 2'd0;
		vns_bankmachine0_state <= 4'd0;
		vns_bankmachine1_state <= 4'd0;
		vns_bankmachine2_state <= 4'd0;
		vns_bankmachine3_state <= 4'd0;
		vns_bankmachine4_state <= 4'd0;
		vns_bankmachine5_state <= 4'd0;
		vns_bankmachine6_state <= 4'd0;
		vns_bankmachine7_state <= 4'd0;
		vns_multiplexer_state <= 4'd0;
		vns_roundrobin0_grant <= 2'd0;
		vns_roundrobin1_grant <= 2'd0;
		vns_roundrobin2_grant <= 2'd0;
		vns_roundrobin3_grant <= 2'd0;
		vns_roundrobin4_grant <= 2'd0;
		vns_roundrobin5_grant <= 2'd0;
		vns_roundrobin6_grant <= 2'd0;
		vns_roundrobin7_grant <= 2'd0;
		vns_rbank <= 3'd0;
		vns_wbank <= 3'd0;
		vns_new_master_wdata_ready0 <= 1'd0;
		vns_new_master_wdata_ready1 <= 1'd0;
		vns_new_master_wdata_ready2 <= 1'd0;
		vns_new_master_wdata_ready3 <= 1'd0;
		vns_new_master_wdata_ready4 <= 1'd0;
		vns_new_master_wdata_ready5 <= 1'd0;
		vns_new_master_wdata_ready6 <= 1'd0;
		vns_new_master_wdata_ready7 <= 1'd0;
		vns_new_master_wdata_ready8 <= 1'd0;
		vns_new_master_rdata_valid0 <= 1'd0;
		vns_new_master_rdata_valid1 <= 1'd0;
		vns_new_master_rdata_valid2 <= 1'd0;
		vns_new_master_rdata_valid3 <= 1'd0;
		vns_new_master_rdata_valid4 <= 1'd0;
		vns_new_master_rdata_valid5 <= 1'd0;
		vns_new_master_rdata_valid6 <= 1'd0;
		vns_new_master_rdata_valid7 <= 1'd0;
		vns_new_master_rdata_valid8 <= 1'd0;
		vns_new_master_rdata_valid9 <= 1'd0;
		vns_new_master_rdata_valid10 <= 1'd0;
		vns_new_master_rdata_valid11 <= 1'd0;
		vns_new_master_rdata_valid12 <= 1'd0;
		vns_new_master_rdata_valid13 <= 1'd0;
		vns_new_master_rdata_valid14 <= 1'd0;
		vns_new_master_rdata_valid15 <= 1'd0;
		vns_new_master_rdata_valid16 <= 1'd0;
		vns_new_master_rdata_valid17 <= 1'd0;
		vns_new_master_rdata_valid18 <= 1'd0;
		vns_new_master_rdata_valid19 <= 1'd0;
		vns_new_master_rdata_valid20 <= 1'd0;
		vns_new_master_rdata_valid21 <= 1'd0;
		vns_new_master_rdata_valid22 <= 1'd0;
		vns_new_master_rdata_valid23 <= 1'd0;
		vns_new_master_rdata_valid24 <= 1'd0;
		vns_new_master_rdata_valid25 <= 1'd0;
		vns_new_master_rdata_valid26 <= 1'd0;
		vns_new_master_rdata_valid27 <= 1'd0;
		vns_new_master_rdata_valid28 <= 1'd0;
		vns_new_master_rdata_valid29 <= 1'd0;
		vns_fullmemorywe_state <= 3'd0;
		vns_litedramwishbone2native_state <= 2'd0;
		vns_edid0_state <= 4'd0;
		vns_edid1_state <= 4'd0;
		vns_dma_state <= 2'd0;
		vns_liteethetherbonepackettx_liteethetherbonepacketpacketizer_state <= 2'd0;
		vns_liteethetherbonepackettx_fsm_state <= 1'd0;
		vns_liteethetherbonepacketrx_liteethetherbonepacketdepacketizer_state <= 2'd0;
		vns_liteethetherbonepacketrx_fsm_state <= 2'd0;
		vns_liteethetherboneprobe_state <= 1'd0;
		vns_liteethetherbonerecorddepacketizer_state <= 1'd0;
		vns_liteethetherbonerecordreceiver_state <= 2'd0;
		vns_liteethetherbonerecordsender_state <= 2'd0;
		vns_liteethetherbonerecordpacketizer_state <= 1'd0;
		vns_liteethetherbonewishbonemaster_state <= 2'd0;
		vns_videooverlaysoc_grant <= 2'd0;
		vns_videooverlaysoc_slave_sel_r <= 5'd0;
		vns_videooverlaysoc_count <= 17'd65536;
		vns_videooverlaysoc_interface0_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface1_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface2_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface3_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_csrbank3_initiator_hres_backstore <= 4'd0;
		vns_videooverlaysoc_csrbank3_initiator_hsync_start_backstore <= 4'd0;
		vns_videooverlaysoc_csrbank3_initiator_hsync_end_backstore <= 4'd0;
		vns_videooverlaysoc_csrbank3_initiator_hscan_backstore <= 4'd0;
		vns_videooverlaysoc_csrbank3_initiator_vres_backstore <= 4'd0;
		vns_videooverlaysoc_csrbank3_initiator_vsync_start_backstore <= 4'd0;
		vns_videooverlaysoc_csrbank3_initiator_vsync_end_backstore <= 4'd0;
		vns_videooverlaysoc_csrbank3_initiator_vscan_backstore <= 4'd0;
		vns_videooverlaysoc_csrbank3_initiator_base_backstore <= 24'd0;
		vns_videooverlaysoc_csrbank3_initiator_length_backstore <= 24'd0;
		vns_videooverlaysoc_sram0_sel_r <= 1'd0;
		vns_videooverlaysoc_interface4_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface5_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_sram1_sel_r <= 1'd0;
		vns_videooverlaysoc_interface6_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface7_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface8_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_sram2_sel_r <= 1'd0;
		vns_videooverlaysoc_interface9_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface10_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface11_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface12_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface13_bank_bus_dat_r <= 8'd0;
		vns_videooverlaysoc_interface14_bank_bus_dat_r <= 8'd0;
	end
	vns_xilinxmultiregimpl0_regs0 <= serial_rx;
	vns_xilinxmultiregimpl0_regs1 <= vns_xilinxmultiregimpl0_regs0;
	vns_xilinxmultiregimpl1_regs0 <= soc_videooverlaysoc_hdmi_in0_freq_q;
	vns_xilinxmultiregimpl1_regs1 <= vns_xilinxmultiregimpl1_regs0;
	vns_xilinxmultiregimpl2_regs0 <= soc_videooverlaysoc_hdmi_in0_edid_hpd_notif_n;
	vns_xilinxmultiregimpl2_regs1 <= vns_xilinxmultiregimpl2_regs0;
	vns_xilinxmultiregimpl3_regs0 <= hdmi_in0_scl;
	vns_xilinxmultiregimpl3_regs1 <= vns_xilinxmultiregimpl3_regs0;
	vns_xilinxmultiregimpl4_regs0 <= soc_videooverlaysoc_hdmi_in0_edid_sda_i_async;
	vns_xilinxmultiregimpl4_regs1 <= vns_xilinxmultiregimpl4_regs0;
	vns_xilinxmultiregimpl5_regs0 <= soc_videooverlaysoc_hdmi_in0_mmcm_locked;
	vns_xilinxmultiregimpl5_regs1 <= vns_xilinxmultiregimpl5_regs0;
	vns_xilinxmultiregimpl11_regs0 <= {soc_videooverlaysoc_hdmi_in0_s7datacapture0_too_early, soc_videooverlaysoc_hdmi_in0_s7datacapture0_too_late};
	vns_xilinxmultiregimpl11_regs1 <= vns_xilinxmultiregimpl11_regs0;
	vns_xilinxmultiregimpl13_regs0 <= soc_videooverlaysoc_hdmi_in0_charsync0_synced;
	vns_xilinxmultiregimpl13_regs1 <= vns_xilinxmultiregimpl13_regs0;
	vns_xilinxmultiregimpl14_regs0 <= soc_videooverlaysoc_hdmi_in0_charsync0_word_sel;
	vns_xilinxmultiregimpl14_regs1 <= vns_xilinxmultiregimpl14_regs0;
	vns_xilinxmultiregimpl15_regs0 <= soc_videooverlaysoc_hdmi_in0_wer0_toggle_i;
	vns_xilinxmultiregimpl15_regs1 <= vns_xilinxmultiregimpl15_regs0;
	vns_xilinxmultiregimpl21_regs0 <= {soc_videooverlaysoc_hdmi_in0_s7datacapture1_too_early, soc_videooverlaysoc_hdmi_in0_s7datacapture1_too_late};
	vns_xilinxmultiregimpl21_regs1 <= vns_xilinxmultiregimpl21_regs0;
	vns_xilinxmultiregimpl23_regs0 <= soc_videooverlaysoc_hdmi_in0_charsync1_synced;
	vns_xilinxmultiregimpl23_regs1 <= vns_xilinxmultiregimpl23_regs0;
	vns_xilinxmultiregimpl24_regs0 <= soc_videooverlaysoc_hdmi_in0_charsync1_word_sel;
	vns_xilinxmultiregimpl24_regs1 <= vns_xilinxmultiregimpl24_regs0;
	vns_xilinxmultiregimpl25_regs0 <= soc_videooverlaysoc_hdmi_in0_wer1_toggle_i;
	vns_xilinxmultiregimpl25_regs1 <= vns_xilinxmultiregimpl25_regs0;
	vns_xilinxmultiregimpl31_regs0 <= {soc_videooverlaysoc_hdmi_in0_s7datacapture2_too_early, soc_videooverlaysoc_hdmi_in0_s7datacapture2_too_late};
	vns_xilinxmultiregimpl31_regs1 <= vns_xilinxmultiregimpl31_regs0;
	vns_xilinxmultiregimpl33_regs0 <= soc_videooverlaysoc_hdmi_in0_charsync2_synced;
	vns_xilinxmultiregimpl33_regs1 <= vns_xilinxmultiregimpl33_regs0;
	vns_xilinxmultiregimpl34_regs0 <= soc_videooverlaysoc_hdmi_in0_charsync2_word_sel;
	vns_xilinxmultiregimpl34_regs1 <= vns_xilinxmultiregimpl34_regs0;
	vns_xilinxmultiregimpl35_regs0 <= soc_videooverlaysoc_hdmi_in0_wer2_toggle_i;
	vns_xilinxmultiregimpl35_regs1 <= vns_xilinxmultiregimpl35_regs0;
	vns_xilinxmultiregimpl36_regs0 <= soc_videooverlaysoc_hdmi_in0_chansync_chan_synced;
	vns_xilinxmultiregimpl36_regs1 <= vns_xilinxmultiregimpl36_regs0;
	vns_xilinxmultiregimpl38_regs0 <= soc_videooverlaysoc_hdmi_in0_resdetection_hcounter_st;
	vns_xilinxmultiregimpl38_regs1 <= vns_xilinxmultiregimpl38_regs0;
	vns_xilinxmultiregimpl39_regs0 <= soc_videooverlaysoc_hdmi_in0_resdetection_vcounter_st;
	vns_xilinxmultiregimpl39_regs1 <= vns_xilinxmultiregimpl39_regs0;
	vns_xilinxmultiregimpl40_regs0 <= soc_videooverlaysoc_hdmi_in1_freq_q;
	vns_xilinxmultiregimpl40_regs1 <= vns_xilinxmultiregimpl40_regs0;
	vns_xilinxmultiregimpl41_regs0 <= (~hdmi_in1_scl);
	vns_xilinxmultiregimpl41_regs1 <= vns_xilinxmultiregimpl41_regs0;
	vns_xilinxmultiregimpl42_regs0 <= soc_videooverlaysoc_hdmi_in1_edid_sda_i_async;
	vns_xilinxmultiregimpl42_regs1 <= vns_xilinxmultiregimpl42_regs0;
	vns_xilinxmultiregimpl43_regs0 <= soc_videooverlaysoc_hdmi_in1_mmcm_locked;
	vns_xilinxmultiregimpl43_regs1 <= vns_xilinxmultiregimpl43_regs0;
	vns_xilinxmultiregimpl49_regs0 <= {soc_videooverlaysoc_hdmi_in1_s7datacapture0_too_early, soc_videooverlaysoc_hdmi_in1_s7datacapture0_too_late};
	vns_xilinxmultiregimpl49_regs1 <= vns_xilinxmultiregimpl49_regs0;
	vns_xilinxmultiregimpl51_regs0 <= soc_videooverlaysoc_hdmi_in1_charsync0_synced;
	vns_xilinxmultiregimpl51_regs1 <= vns_xilinxmultiregimpl51_regs0;
	vns_xilinxmultiregimpl52_regs0 <= soc_videooverlaysoc_hdmi_in1_charsync0_word_sel;
	vns_xilinxmultiregimpl52_regs1 <= vns_xilinxmultiregimpl52_regs0;
	vns_xilinxmultiregimpl53_regs0 <= soc_videooverlaysoc_hdmi_in1_wer0_toggle_i;
	vns_xilinxmultiregimpl53_regs1 <= vns_xilinxmultiregimpl53_regs0;
	vns_xilinxmultiregimpl59_regs0 <= {soc_videooverlaysoc_hdmi_in1_s7datacapture1_too_early, soc_videooverlaysoc_hdmi_in1_s7datacapture1_too_late};
	vns_xilinxmultiregimpl59_regs1 <= vns_xilinxmultiregimpl59_regs0;
	vns_xilinxmultiregimpl61_regs0 <= soc_videooverlaysoc_hdmi_in1_charsync1_synced;
	vns_xilinxmultiregimpl61_regs1 <= vns_xilinxmultiregimpl61_regs0;
	vns_xilinxmultiregimpl62_regs0 <= soc_videooverlaysoc_hdmi_in1_charsync1_word_sel;
	vns_xilinxmultiregimpl62_regs1 <= vns_xilinxmultiregimpl62_regs0;
	vns_xilinxmultiregimpl63_regs0 <= soc_videooverlaysoc_hdmi_in1_wer1_toggle_i;
	vns_xilinxmultiregimpl63_regs1 <= vns_xilinxmultiregimpl63_regs0;
	vns_xilinxmultiregimpl69_regs0 <= {soc_videooverlaysoc_hdmi_in1_s7datacapture2_too_early, soc_videooverlaysoc_hdmi_in1_s7datacapture2_too_late};
	vns_xilinxmultiregimpl69_regs1 <= vns_xilinxmultiregimpl69_regs0;
	vns_xilinxmultiregimpl71_regs0 <= soc_videooverlaysoc_hdmi_in1_charsync2_synced;
	vns_xilinxmultiregimpl71_regs1 <= vns_xilinxmultiregimpl71_regs0;
	vns_xilinxmultiregimpl72_regs0 <= soc_videooverlaysoc_hdmi_in1_charsync2_word_sel;
	vns_xilinxmultiregimpl72_regs1 <= vns_xilinxmultiregimpl72_regs0;
	vns_xilinxmultiregimpl73_regs0 <= soc_videooverlaysoc_hdmi_in1_wer2_toggle_i;
	vns_xilinxmultiregimpl73_regs1 <= vns_xilinxmultiregimpl73_regs0;
	vns_xilinxmultiregimpl74_regs0 <= soc_videooverlaysoc_hdmi_in1_chansync_chan_synced;
	vns_xilinxmultiregimpl74_regs1 <= vns_xilinxmultiregimpl74_regs0;
	vns_xilinxmultiregimpl76_regs0 <= soc_videooverlaysoc_hdmi_in1_resdetection_hcounter_st;
	vns_xilinxmultiregimpl76_regs1 <= vns_xilinxmultiregimpl76_regs0;
	vns_xilinxmultiregimpl77_regs0 <= soc_videooverlaysoc_hdmi_in1_resdetection_vcounter_st;
	vns_xilinxmultiregimpl77_regs1 <= vns_xilinxmultiregimpl77_regs0;
	vns_xilinxmultiregimpl78_regs0 <= soc_videooverlaysoc_hdmi_in1_frame_graycounter0_q;
	vns_xilinxmultiregimpl78_regs1 <= vns_xilinxmultiregimpl78_regs0;
	vns_xilinxmultiregimpl80_regs0 <= soc_videooverlaysoc_hdmi_in1_frame_pix_overflow;
	vns_xilinxmultiregimpl80_regs1 <= vns_xilinxmultiregimpl80_regs0;
	vns_xilinxmultiregimpl82_regs0 <= soc_videooverlaysoc_hdmi_in1_frame_overflow_reset_ack_toggle_i;
	vns_xilinxmultiregimpl82_regs1 <= vns_xilinxmultiregimpl82_regs0;
	vns_xilinxmultiregimpl83_regs0 <= soc_videooverlaysoc_out_dram_port_cmd_fifo_graycounter0_q;
	vns_xilinxmultiregimpl83_regs1 <= vns_xilinxmultiregimpl83_regs0;
	vns_xilinxmultiregimpl86_regs0 <= soc_videooverlaysoc_out_dram_port_rdata_fifo_graycounter1_q;
	vns_xilinxmultiregimpl86_regs1 <= vns_xilinxmultiregimpl86_regs0;
	vns_xilinxmultiregimpl88_regs0 <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_graycounter1_q;
	vns_xilinxmultiregimpl88_regs1 <= vns_xilinxmultiregimpl88_regs0;
	vns_xilinxmultiregimpl89_regs0 <= soc_videooverlaysoc_hdmi_core_out0_underflow_enable_storage;
	vns_xilinxmultiregimpl89_regs1 <= vns_xilinxmultiregimpl89_regs0;
end

VexRiscv VexRiscv(
	.clk(sys_clk),
	.dBusWishbone_ACK(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_ack),
	.dBusWishbone_DAT_MISO(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_dat_r),
	.dBusWishbone_ERR(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_d_err),
	.debugReset(sys_rst),
	.debug_bus_cmd_payload_address(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_address),
	.debug_bus_cmd_payload_data(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_data),
	.debug_bus_cmd_payload_wr(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_payload_wr),
	.debug_bus_cmd_valid(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_cmd_valid),
	.externalInterruptArray(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_interrupt),
	.externalResetVector(1'd0),
	.iBusWishbone_ACK(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_ack),
	.iBusWishbone_DAT_MISO(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_dat_r),
	.iBusWishbone_ERR(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_i_err),
	.reset((soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_cpu_reset | soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_reset)),
	.timerInterrupt(1'd0),
	.dBusWishbone_ADR(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_adr),
	.dBusWishbone_BTE(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_bte),
	.dBusWishbone_CTI(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_cti),
	.dBusWishbone_CYC(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_cyc),
	.dBusWishbone_DAT_MOSI(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_dat_w),
	.dBusWishbone_SEL(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_sel),
	.dBusWishbone_STB(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_stb),
	.dBusWishbone_WE(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_dbus_we),
	.debug_bus_cmd_ready(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_o_cmd_ready),
	.debug_bus_rsp_data(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_o_rsp_data),
	.debug_resetOut(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_o_resetOut),
	.iBusWishbone_ADR(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_adr),
	.iBusWishbone_BTE(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_bte),
	.iBusWishbone_CTI(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_cti),
	.iBusWishbone_CYC(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_cyc),
	.iBusWishbone_DAT_MOSI(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_dat_w),
	.iBusWishbone_SEL(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_sel),
	.iBusWishbone_STB(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_stb),
	.iBusWishbone_WE(soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_vexriscv_ibus_we)
);

reg [31:0] mem[0:5119];
reg [12:0] memadr;
always @(posedge sys_clk) begin
	memadr <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_rom_dat_r = mem[memadr];

initial begin
	$readmemh("mem.init", mem);
end

reg [31:0] mem_1[0:4095];
reg [11:0] memadr_1;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_we[0])
		mem_1[soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_adr][7:0] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_dat_w[7:0];
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_we[1])
		mem_1[soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_adr][15:8] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_dat_w[15:8];
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_we[2])
		mem_1[soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_adr][23:16] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_dat_w[23:16];
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_we[3])
		mem_1[soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_adr][31:24] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_dat_w[31:24];
	memadr_1 <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_sram_dat_r = mem_1[memadr_1];

reg [9:0] storage[0:15];
reg [9:0] memdat;
reg [9:0] memdat_1;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_we)
		storage[soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_adr] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_dat_w;
	memdat <= storage[soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_rdport_re)
		memdat_1 <= storage[soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_rdport_adr];
end

assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_wrport_dat_r = memdat;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_tx_fifo_rdport_dat_r = memdat_1;

reg [9:0] storage_1[0:15];
reg [9:0] memdat_2;
reg [9:0] memdat_3;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_we)
		storage_1[soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_adr] <= soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_dat_w;
	memdat_2 <= storage_1[soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_rdport_re)
		memdat_3 <= storage_1[soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_rdport_adr];
end

assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_wrport_dat_r = memdat_2;
assign soc_videooverlaysoc_videooverlaysoc_videooverlaysoc_uart_rx_fifo_rdport_dat_r = memdat_3;

reg [7:0] mem_2[0:20];
reg [4:0] memadr_2;
always @(posedge sys_clk) begin
	memadr_2 <= vns_videooverlaysoc_sram2_adr;
end

assign vns_videooverlaysoc_sram2_dat_r = mem_2[memadr_2];

initial begin
	$readmemh("mem_2.init", mem_2);
end

PLLE2_BASE #(
	.CLKFBOUT_MULT(6'd32),
	.CLKIN1_PERIOD(20.0),
	.CLKOUT0_DIVIDE(5'd16),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(3'd4),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(3'd4),
	.CLKOUT2_PHASE(90.0),
	.CLKOUT3_DIVIDE(4'd8),
	.CLKOUT3_PHASE(0.0),
	.CLKOUT4_DIVIDE(6'd32),
	.CLKOUT4_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01),
	.STARTUP_WAIT("FALSE")
) PLLE2_BASE (
	.CLKFBIN(soc_videooverlaysoc_videooverlaysoc_crg_pll_fb_bufg),
	.CLKIN1(clk50),
	.CLKFBOUT(soc_videooverlaysoc_videooverlaysoc_crg_pll_fb),
	.CLKOUT0(soc_videooverlaysoc_videooverlaysoc_crg_pll_sys),
	.CLKOUT1(soc_videooverlaysoc_videooverlaysoc_crg_pll_sys4x),
	.CLKOUT2(soc_videooverlaysoc_videooverlaysoc_crg_pll_sys4x_dqs),
	.CLKOUT3(soc_videooverlaysoc_videooverlaysoc_crg_pll_clk200),
	.CLKOUT4(soc_videooverlaysoc_videooverlaysoc_crg_pll_clk50),
	.LOCKED(soc_videooverlaysoc_videooverlaysoc_crg_pll_locked)
);

BUFG BUFG(
	.I(soc_videooverlaysoc_videooverlaysoc_crg_pll_sys),
	.O(sys_clk)
);

BUFG BUFG_1(
	.I(soc_videooverlaysoc_videooverlaysoc_crg_pll_fb),
	.O(soc_videooverlaysoc_videooverlaysoc_crg_pll_fb_bufg)
);

BUFG BUFG_2(
	.I(soc_videooverlaysoc_videooverlaysoc_crg_pll_clk200),
	.O(clk200_clk)
);

BUFG BUFG_3(
	.I(soc_videooverlaysoc_videooverlaysoc_crg_pll_sys4x),
	.O(sys4x_clk)
);

BUFG BUFG_4(
	.I(soc_videooverlaysoc_videooverlaysoc_crg_pll_sys4x_dqs),
	.O(sys4x_dqs_clk)
);

BUFG BUFG_5(
	.I(soc_videooverlaysoc_videooverlaysoc_crg_pll_clk50),
	.O(eth_clk)
);

IDELAYCTRL IDELAYCTRL(
	.REFCLK(clk200_clk),
	.RST(soc_videooverlaysoc_videooverlaysoc_crg_ic_reset)
);

XADC #(
	.INIT_40(16'd36864),
	.INIT_41(14'd12016),
	.INIT_42(11'd1024),
	.INIT_48(15'd18177),
	.INIT_49(4'd15),
	.INIT_4A(15'd18176),
	.INIT_4B(1'd0),
	.INIT_4C(1'd0),
	.INIT_4D(1'd0),
	.INIT_4E(1'd0),
	.INIT_4F(1'd0),
	.INIT_50(16'd46573),
	.INIT_51(15'd22937),
	.INIT_52(16'd41287),
	.INIT_53(16'd56797),
	.INIT_54(16'd43322),
	.INIT_55(15'd20753),
	.INIT_56(16'd37355),
	.INIT_57(16'd44622),
	.INIT_58(15'd22937),
	.INIT_5C(15'd20753)
) XADC (
	.CONVST(1'd0),
	.CONVSTCLK(1'd0),
	.DADDR(soc_videooverlaysoc_videooverlaysoc_channel),
	.DCLK(sys_clk),
	.DEN(soc_videooverlaysoc_videooverlaysoc_eoc),
	.DI(1'd0),
	.DWE(1'd0),
	.RESET(sys_rst),
	.VAUXN(1'd0),
	.VAUXP(1'd1),
	.VN(1'd0),
	.VP(1'd1),
	.ALM(soc_videooverlaysoc_videooverlaysoc_alarm),
	.BUSY(soc_videooverlaysoc_videooverlaysoc_busy),
	.CHANNEL(soc_videooverlaysoc_videooverlaysoc_channel),
	.DO(soc_videooverlaysoc_videooverlaysoc_data),
	.DRDY(soc_videooverlaysoc_videooverlaysoc_drdy),
	.EOC(soc_videooverlaysoc_videooverlaysoc_eoc),
	.EOS(soc_videooverlaysoc_videooverlaysoc_eos),
	.OT(soc_videooverlaysoc_videooverlaysoc_ot)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(1'd0),
	.D2(1'd1),
	.D3(1'd0),
	.D4(1'd1),
	.D5(1'd0),
	.D6(1'd1),
	.D7(1'd0),
	.D8(1'd1),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_sd_clk_se)
);

OBUFDS OBUFDS(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_sd_clk_se),
	.O(ddram_clk_p),
	.OB(ddram_clk_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_1 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[0]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[0]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[0]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[0]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[0]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[0]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[0]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[1]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[1]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[1]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[1]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[1]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[1]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[1]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_3 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[2]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[2]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[2]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[2]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[2]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[2]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[2]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_4 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[3]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[3]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[3]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[3]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[3]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[3]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[3]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[3])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_5 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[4]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[4]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[4]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[4]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[4]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[4]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[4]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[4]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[4])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_6 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[5]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[5]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[5]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[5]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[5]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[5]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[5]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[5]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[5])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_7 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[6]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[6]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[6]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[6]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[6]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[6]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[6]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[6]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[6])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_8 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[7]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[7]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[7]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[7]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[7]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[7]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[7]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[7])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_9 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[8]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[8]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[8]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[8]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[8]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[8]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[8]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[8]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[8])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_10 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[9]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[9]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[9]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[9]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[9]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[9]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[9]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[9]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[9])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_11 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[10]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[10]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[10]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[10]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[10]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[10]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[10]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[10]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[10])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_12 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[11]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[11]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[11]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[11]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[11]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[11]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[11]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[11]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[11])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_13 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[12]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[12]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[12]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[12]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[12]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[12]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[12]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[12]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[12])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_14 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[13]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_address[13]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[13]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_address[13]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[13]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_address[13]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[13]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_address[13]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[13])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_15 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_bank[0]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_bank[0]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_bank[0]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_bank[0]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_bank[0]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_bank[0]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_bank[0]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_bank[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_16 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_bank[1]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_bank[1]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_bank[1]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_bank[1]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_bank[1]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_bank[1]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_bank[1]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_bank[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_17 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_bank[2]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_bank[2]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_bank[2]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_bank[2]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_bank[2]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_bank[2]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_bank[2]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_bank[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_18 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_ras_n),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_ras_n),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_ras_n),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_ras_n),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_ras_n),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_ras_n),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_ras_n),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_ras_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ras_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_19 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cas_n),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cas_n),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cas_n),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cas_n),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cas_n),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cas_n),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cas_n),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cas_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cas_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_20 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_we_n),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_we_n),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_we_n),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_we_n),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_we_n),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_we_n),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_we_n),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_we_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_we_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_21 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cke),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cke),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cke),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cke),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cke),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cke),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cke),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cke),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cke)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_22 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_odt),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_odt),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_odt),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_odt),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_odt),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_odt),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_odt),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_odt),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_odt)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_23 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_reset_n),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_reset_n),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_reset_n),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_reset_n),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_reset_n),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_reset_n),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_reset_n),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_reset_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_reset_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_24 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cs_n),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_cs_n),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cs_n),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_cs_n),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cs_n),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_cs_n),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cs_n),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_cs_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cs_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_25 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_mask[0]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_mask[4]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_mask[0]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_mask[4]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_mask[0]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_mask[4]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_mask[0]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_mask[4]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_26 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[0]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[1]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[2]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[3]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[4]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[5]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[6]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(soc_videooverlaysoc_videooverlaysoc_a7ddrphy0),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay0),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t0)
);

OBUFTDS OBUFTDS(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay0),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t0),
	.O(ddram_dqs_p[0]),
	.OB(ddram_dqs_n[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_27 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_mask[1]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_mask[5]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_mask[1]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_mask[5]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_mask[1]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_mask[5]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_mask[1]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_mask[5]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_28 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[0]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[1]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[2]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[3]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[4]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[5]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[6]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(soc_videooverlaysoc_videooverlaysoc_a7ddrphy1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay1),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t1)
);

OBUFTDS OBUFTDS_1(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay1),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t1),
	.O(ddram_dqs_p[1]),
	.OB(ddram_dqs_n[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_29 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_mask[2]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_mask[6]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_mask[2]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_mask[6]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_mask[2]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_mask[6]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_mask[2]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_mask[6]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_30 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[0]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[1]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[2]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[3]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[4]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[5]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[6]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(soc_videooverlaysoc_videooverlaysoc_a7ddrphy2),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay2),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t2)
);

OBUFTDS OBUFTDS_2(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay2),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t2),
	.O(ddram_dqs_p[2]),
	.OB(ddram_dqs_n[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_31 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_mask[3]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata_mask[7]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_mask[3]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata_mask[7]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_mask[3]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata_mask[7]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_mask[3]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata_mask[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[3])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_32 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[0]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[1]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[2]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[3]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[4]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[5]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[6]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(soc_videooverlaysoc_videooverlaysoc_a7ddrphy3),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay3),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t3)
);

OBUFTDS OBUFTDS_3(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_nodelay3),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dqs_t3),
	.O(ddram_dqs_p[3]),
	.OB(ddram_dqs_n[3])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_33 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[0]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[32]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[0]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[32]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[0]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[32]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[0]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[32]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay0),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed0),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data0[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data0[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data0[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data0[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data0[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data0[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data0[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data0[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay0),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed0)
);

IOBUF IOBUF(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay0),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t0),
	.IO(ddram_dq[0]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_34 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[1]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[33]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[1]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[33]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[1]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[33]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[1]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[33]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay1),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t1)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_1 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed1),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data1[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data1[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data1[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data1[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data1[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data1[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data1[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data1[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_1 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay1),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed1)
);

IOBUF IOBUF_1(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay1),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t1),
	.IO(ddram_dq[1]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_35 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[2]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[34]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[2]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[34]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[2]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[34]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[2]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[34]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay2),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t2)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_2 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed2),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data2[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data2[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data2[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data2[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data2[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data2[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data2[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data2[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_2 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay2),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed2)
);

IOBUF IOBUF_2(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay2),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t2),
	.IO(ddram_dq[2]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_36 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[3]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[35]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[3]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[35]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[3]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[35]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[3]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[35]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay3),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t3)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_3 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed3),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data3[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data3[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data3[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data3[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data3[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data3[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data3[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data3[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_3 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay3),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed3)
);

IOBUF IOBUF_3(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay3),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t3),
	.IO(ddram_dq[3]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_37 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[4]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[36]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[4]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[36]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[4]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[36]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[4]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[36]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay4),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t4)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_4 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed4),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data4[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data4[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data4[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data4[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data4[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data4[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data4[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data4[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_4 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay4),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed4)
);

IOBUF IOBUF_4(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay4),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t4),
	.IO(ddram_dq[4]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_38 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[5]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[37]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[5]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[37]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[5]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[37]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[5]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[37]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay5),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t5)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_5 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed5),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data5[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data5[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data5[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data5[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data5[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data5[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data5[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data5[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_5 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay5),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed5)
);

IOBUF IOBUF_5(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay5),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t5),
	.IO(ddram_dq[5]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_39 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[6]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[38]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[6]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[38]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[6]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[38]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[6]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[38]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay6),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t6)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_6 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed6),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data6[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data6[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data6[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data6[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data6[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data6[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data6[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data6[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_6 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay6),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed6)
);

IOBUF IOBUF_6(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay6),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t6),
	.IO(ddram_dq[6]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_40 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[7]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[39]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[7]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[39]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[7]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[39]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[7]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[39]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay7),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t7)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_7 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed7),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data7[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data7[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data7[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data7[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data7[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data7[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data7[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data7[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_7 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay7),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[0] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed7)
);

IOBUF IOBUF_7(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay7),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t7),
	.IO(ddram_dq[7]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay7)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_41 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[8]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[40]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[8]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[40]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[8]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[40]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[8]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[40]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay8),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t8)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_8 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed8),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data8[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data8[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data8[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data8[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data8[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data8[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data8[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data8[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_8 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay8),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed8)
);

IOBUF IOBUF_8(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay8),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t8),
	.IO(ddram_dq[8]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay8)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_42 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[9]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[41]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[9]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[41]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[9]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[41]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[9]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[41]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay9),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t9)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_9 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed9),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data9[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data9[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data9[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data9[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data9[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data9[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data9[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data9[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_9 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay9),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed9)
);

IOBUF IOBUF_9(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay9),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t9),
	.IO(ddram_dq[9]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay9)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_43 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[10]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[42]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[10]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[42]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[10]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[42]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[10]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[42]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay10),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t10)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_10 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed10),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data10[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data10[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data10[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data10[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data10[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data10[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data10[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data10[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_10 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay10),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed10)
);

IOBUF IOBUF_10(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay10),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t10),
	.IO(ddram_dq[10]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay10)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_44 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[11]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[43]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[11]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[43]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[11]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[43]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[11]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[43]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay11),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t11)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_11 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed11),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data11[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data11[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data11[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data11[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data11[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data11[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data11[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data11[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_11 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay11),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed11)
);

IOBUF IOBUF_11(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay11),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t11),
	.IO(ddram_dq[11]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay11)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_45 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[12]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[44]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[12]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[44]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[12]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[44]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[12]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[44]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay12),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t12)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_12 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed12),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data12[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data12[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data12[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data12[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data12[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data12[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data12[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data12[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_12 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay12),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed12)
);

IOBUF IOBUF_12(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay12),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t12),
	.IO(ddram_dq[12]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay12)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_46 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[13]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[45]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[13]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[45]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[13]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[45]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[13]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[45]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay13),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t13)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_13 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed13),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data13[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data13[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data13[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data13[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data13[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data13[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data13[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data13[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_13 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay13),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed13)
);

IOBUF IOBUF_13(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay13),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t13),
	.IO(ddram_dq[13]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay13)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_47 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[14]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[46]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[14]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[46]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[14]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[46]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[14]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[46]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay14),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t14)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_14 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed14),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data14[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data14[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data14[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data14[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data14[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data14[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data14[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data14[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_14 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay14),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed14)
);

IOBUF IOBUF_14(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay14),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t14),
	.IO(ddram_dq[14]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay14)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_48 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[15]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[47]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[15]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[47]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[15]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[47]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[15]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[47]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay15),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t15)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_15 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed15),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data15[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data15[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data15[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data15[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data15[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data15[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data15[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data15[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_15 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay15),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[1] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed15)
);

IOBUF IOBUF_15(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay15),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t15),
	.IO(ddram_dq[15]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay15)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_49 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[16]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[48]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[16]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[48]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[16]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[48]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[16]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[48]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay16),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t16)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_16 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed16),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data16[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data16[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data16[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data16[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data16[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data16[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data16[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data16[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_16 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay16),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed16)
);

IOBUF IOBUF_16(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay16),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t16),
	.IO(ddram_dq[16]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay16)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_50 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[17]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[49]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[17]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[49]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[17]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[49]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[17]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[49]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay17),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t17)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_17 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed17),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data17[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data17[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data17[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data17[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data17[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data17[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data17[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data17[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_17 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay17),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed17)
);

IOBUF IOBUF_17(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay17),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t17),
	.IO(ddram_dq[17]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay17)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_51 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[18]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[50]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[18]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[50]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[18]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[50]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[18]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[50]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay18),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t18)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_18 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed18),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data18[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data18[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data18[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data18[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data18[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data18[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data18[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data18[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_18 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay18),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed18)
);

IOBUF IOBUF_18(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay18),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t18),
	.IO(ddram_dq[18]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay18)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_52 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[19]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[51]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[19]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[51]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[19]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[51]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[19]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[51]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay19),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t19)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_19 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed19),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data19[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data19[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data19[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data19[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data19[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data19[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data19[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data19[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_19 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay19),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed19)
);

IOBUF IOBUF_19(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay19),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t19),
	.IO(ddram_dq[19]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay19)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_53 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[20]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[52]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[20]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[52]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[20]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[52]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[20]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[52]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay20),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t20)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_20 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed20),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data20[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data20[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data20[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data20[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data20[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data20[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data20[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data20[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_20 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay20),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed20)
);

IOBUF IOBUF_20(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay20),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t20),
	.IO(ddram_dq[20]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay20)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_54 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[21]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[53]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[21]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[53]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[21]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[53]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[21]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[53]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay21),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t21)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_21 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed21),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data21[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data21[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data21[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data21[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data21[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data21[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data21[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data21[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_21 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay21),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed21)
);

IOBUF IOBUF_21(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay21),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t21),
	.IO(ddram_dq[21]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay21)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_55 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[22]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[54]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[22]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[54]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[22]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[54]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[22]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[54]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay22),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t22)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_22 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed22),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data22[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data22[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data22[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data22[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data22[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data22[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data22[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data22[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_22 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay22),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed22)
);

IOBUF IOBUF_22(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay22),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t22),
	.IO(ddram_dq[22]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay22)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_56 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[23]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[55]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[23]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[55]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[23]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[55]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[23]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[55]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay23),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t23)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_23 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed23),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data23[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data23[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data23[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data23[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data23[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data23[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data23[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data23[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_23 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay23),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[2] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed23)
);

IOBUF IOBUF_23(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay23),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t23),
	.IO(ddram_dq[23]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay23)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_57 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[24]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[56]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[24]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[56]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[24]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[56]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[24]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[56]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay24),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t24)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_24 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed24),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data24[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data24[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data24[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data24[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data24[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data24[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data24[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data24[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_24 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay24),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed24)
);

IOBUF IOBUF_24(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay24),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t24),
	.IO(ddram_dq[24]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay24)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_58 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[25]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[57]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[25]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[57]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[25]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[57]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[25]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[57]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay25),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t25)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_25 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed25),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data25[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data25[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data25[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data25[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data25[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data25[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data25[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data25[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_25 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay25),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed25)
);

IOBUF IOBUF_25(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay25),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t25),
	.IO(ddram_dq[25]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay25)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_59 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[26]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[58]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[26]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[58]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[26]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[58]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[26]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[58]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay26),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t26)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_26 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed26),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data26[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data26[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data26[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data26[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data26[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data26[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data26[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data26[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_26 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay26),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed26)
);

IOBUF IOBUF_26(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay26),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t26),
	.IO(ddram_dq[26]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay26)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_60 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[27]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[59]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[27]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[59]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[27]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[59]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[27]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[59]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay27),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t27)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_27 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed27),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data27[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data27[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data27[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data27[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data27[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data27[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data27[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data27[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_27 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay27),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed27)
);

IOBUF IOBUF_27(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay27),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t27),
	.IO(ddram_dq[27]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay27)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_61 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[28]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[60]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[28]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[60]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[28]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[60]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[28]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[60]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay28),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t28)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_28 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed28),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data28[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data28[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data28[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data28[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data28[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data28[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data28[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data28[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_28 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay28),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed28)
);

IOBUF IOBUF_28(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay28),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t28),
	.IO(ddram_dq[28]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay28)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_62 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[29]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[61]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[29]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[61]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[29]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[61]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[29]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[61]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay29),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t29)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_29 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed29),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data29[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data29[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data29[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data29[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data29[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data29[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data29[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data29[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_29 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay29),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed29)
);

IOBUF IOBUF_29(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay29),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t29),
	.IO(ddram_dq[29]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay29)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_63 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[30]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[62]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[30]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[62]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[30]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[62]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[30]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[62]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay30),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t30)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_30 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed30),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data30[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data30[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data30[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data30[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data30[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data30[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data30[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data30[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_30 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay30),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed30)
);

IOBUF IOBUF_30(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay30),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t30),
	.IO(ddram_dq[30]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay30)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_64 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[31]),
	.D2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p0_wrdata[63]),
	.D3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[31]),
	.D4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p1_wrdata[63]),
	.D5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[31]),
	.D6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p2_wrdata[63]),
	.D7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[31]),
	.D8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dfi_p3_wrdata[63]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videooverlaysoc_videooverlaysoc_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay31),
	.TQ(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t31)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_31 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed31),
	.RST(sys_rst),
	.Q1(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data31[7]),
	.Q2(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data31[6]),
	.Q3(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data31[5]),
	.Q4(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data31[4]),
	.Q5(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data31[3]),
	.Q6(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data31[2]),
	.Q7(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data31[1]),
	.Q8(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_data31[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_31 (
	.C(sys_clk),
	.CE((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay31),
	.INC(1'd1),
	.LD((soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dly_sel_storage[3] & soc_videooverlaysoc_videooverlaysoc_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_delayed31)
);

IOBUF IOBUF_31(
	.I(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_o_nodelay31),
	.T(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_t31),
	.IO(ddram_dq[31]),
	.O(soc_videooverlaysoc_videooverlaysoc_a7ddrphy_dq_i_nodelay31)
);

reg [23:0] storage_2[0:7];
reg [23:0] memdat_4;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_we)
		storage_2[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr] <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_dat_w;
	memdat_4 <= storage_2[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_wrport_dat_r = memdat_4;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_rdport_dat_r = storage_2[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine0_cmd_buffer_lookahead_rdport_adr];

reg [23:0] storage_3[0:7];
reg [23:0] memdat_5;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_we)
		storage_3[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr] <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_dat_w;
	memdat_5 <= storage_3[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_wrport_dat_r = memdat_5;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_rdport_dat_r = storage_3[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine1_cmd_buffer_lookahead_rdport_adr];

reg [23:0] storage_4[0:7];
reg [23:0] memdat_6;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_we)
		storage_4[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr] <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_dat_w;
	memdat_6 <= storage_4[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_wrport_dat_r = memdat_6;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_rdport_dat_r = storage_4[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine2_cmd_buffer_lookahead_rdport_adr];

reg [23:0] storage_5[0:7];
reg [23:0] memdat_7;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_we)
		storage_5[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr] <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_dat_w;
	memdat_7 <= storage_5[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_wrport_dat_r = memdat_7;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_rdport_dat_r = storage_5[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine3_cmd_buffer_lookahead_rdport_adr];

reg [23:0] storage_6[0:7];
reg [23:0] memdat_8;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_we)
		storage_6[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr] <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_dat_w;
	memdat_8 <= storage_6[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_wrport_dat_r = memdat_8;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_rdport_dat_r = storage_6[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine4_cmd_buffer_lookahead_rdport_adr];

reg [23:0] storage_7[0:7];
reg [23:0] memdat_9;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_we)
		storage_7[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr] <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_dat_w;
	memdat_9 <= storage_7[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_wrport_dat_r = memdat_9;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_rdport_dat_r = storage_7[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine5_cmd_buffer_lookahead_rdport_adr];

reg [23:0] storage_8[0:7];
reg [23:0] memdat_10;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_we)
		storage_8[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr] <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_dat_w;
	memdat_10 <= storage_8[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_wrport_dat_r = memdat_10;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_rdport_dat_r = storage_8[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine6_cmd_buffer_lookahead_rdport_adr];

reg [23:0] storage_9[0:7];
reg [23:0] memdat_11;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_we)
		storage_9[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr] <= soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_dat_w;
	memdat_11 <= storage_9[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_wrport_dat_r = memdat_11;
assign soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_rdport_dat_r = storage_9[soc_videooverlaysoc_videooverlaysoc_sdram_bankmachine7_cmd_buffer_lookahead_rdport_adr];

reg [25:0] tag_mem[0:255];
reg [7:0] memadr_3;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_tag_port_we)
		tag_mem[soc_videooverlaysoc_videooverlaysoc_tag_port_adr] <= soc_videooverlaysoc_videooverlaysoc_tag_port_dat_w;
	memadr_3 <= soc_videooverlaysoc_videooverlaysoc_tag_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_tag_port_dat_r = tag_mem[memadr_3];

reg [7:0] edid_mem[0:255];
reg [7:0] memadr_4;
reg [7:0] memadr_5;
always @(posedge sys_clk) begin
	memadr_4 <= soc_videooverlaysoc_hdmi_in0_edid_adr;
end

always @(posedge sys_clk) begin
	if (vns_videooverlaysoc_sram0_we)
		edid_mem[vns_videooverlaysoc_sram0_adr] <= vns_videooverlaysoc_sram0_dat_w;
	memadr_5 <= vns_videooverlaysoc_sram0_adr;
end

assign soc_videooverlaysoc_hdmi_in0_edid_dat_r = edid_mem[memadr_4];
assign vns_videooverlaysoc_sram0_dat_r = edid_mem[memadr_5];

initial begin
	$readmemh("edid_mem.init", edid_mem);
end

assign hdmi_in0_sda = soc_videooverlaysoc_hdmi_in0_edid_sda_drv_reg ? 1'd0 : 1'bz;
assign soc_videooverlaysoc_hdmi_in0_edid_sda_i_async = hdmi_in0_sda;

IBUFDS_DIFF_OUT hdmi_in_ibufds(
	.I(hdmi_in0_clk_p),
	.IB(hdmi_in0_clk_n),
	.OB(soc_videooverlaysoc_hdmi_in0_clk_input)
);

BUFR BUFR(
	.I(soc_videooverlaysoc_hdmi_in0_clk_input),
	.O(soc_videooverlaysoc_hdmi_in0_clk_input_bufr)
);

MMCME2_ADV #(
	.BANDWIDTH("OPTIMIZED"),
	.CLKFBOUT_MULT_F(5.0),
	.CLKFBOUT_PHASE(0.0),
	.CLKIN1_PERIOD(6.734),
	.CLKOUT0_DIVIDE_F(3'd5),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(3'd4),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(1'd1),
	.CLKOUT2_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01)
) MMCME2_ADV (
	.CLKFBIN(soc_videooverlaysoc_hdmi_in0_mmcm_fb_o),
	.CLKIN1(soc_videooverlaysoc_hdmi_in0_clk_input_bufr),
	.DADDR(soc_videooverlaysoc_hdmi_in0_mmcm_adr_storage),
	.DCLK(sys_clk),
	.DEN((soc_videooverlaysoc_hdmi_in0_mmcm_read_re | soc_videooverlaysoc_hdmi_in0_mmcm_write_re)),
	.DI(soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage),
	.DWE(soc_videooverlaysoc_hdmi_in0_mmcm_write_re),
	.RST(soc_videooverlaysoc_hdmi_in0_mmcm_reset_storage),
	.CLKFBOUT(soc_videooverlaysoc_hdmi_in0_mmcm_fb),
	.CLKOUT0(soc_videooverlaysoc_hdmi_in0_mmcm_clk0),
	.CLKOUT1(soc_videooverlaysoc_hdmi_in0_mmcm_clk1),
	.CLKOUT2(soc_videooverlaysoc_hdmi_in0_mmcm_clk2),
	.DO(soc_videooverlaysoc_hdmi_in0_mmcm_dat_r_status),
	.DRDY(soc_videooverlaysoc_hdmi_in0_mmcm_drdy),
	.LOCKED(soc_videooverlaysoc_hdmi_in0_mmcm_locked)
);

BUFG BUFG_6(
	.I(soc_videooverlaysoc_hdmi_in0_mmcm_clk0),
	.O(hdmi_in0_pix_clk)
);

BUFG BUFG_7(
	.I(soc_videooverlaysoc_hdmi_in0_mmcm_clk1),
	.O(hdmi_in0_pix1p25x_clk)
);

BUFIO BUFIO(
	.I(soc_videooverlaysoc_hdmi_in0_mmcm_clk2),
	.O(hdmi_in0_pix5x_clk)
);

BUFG BUFG_8(
	.I(soc_videooverlaysoc_hdmi_in0_mmcm_fb),
	.O(soc_videooverlaysoc_hdmi_in0_mmcm_fb_o)
);

PLLE2_ADV #(
	.BANDWIDTH("LOW"),
	.CLKFBOUT_MULT(4'd10),
	.CLKFBOUT_PHASE(0.0),
	.CLKIN1_PERIOD(6.734),
	.CLKOUT0_DIVIDE(4'd10),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT2_DIVIDE(2'd2),
	.CLKOUT2_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01)
) PLLE2_ADV (
	.CLKFBIN(soc_videooverlaysoc_hdmi_in0_mmcm_fb2_o),
	.CLKIN1(soc_videooverlaysoc_hdmi_in0_mmcm_clk0),
	.DADDR(soc_videooverlaysoc_hdmi_in0_mmcm_adr_storage),
	.DCLK(sys_clk),
	.DEN((soc_videooverlaysoc_hdmi_in0_mmcm_read_o_re | soc_videooverlaysoc_hdmi_in0_mmcm_write_o_re)),
	.DI(soc_videooverlaysoc_hdmi_in0_mmcm_dat_w_storage),
	.DWE(soc_videooverlaysoc_hdmi_in0_mmcm_write_o_re),
	.RST(soc_videooverlaysoc_hdmi_in0_mmcm_reset_storage),
	.CLKFBOUT(soc_videooverlaysoc_hdmi_in0_mmcm_fb2_o),
	.CLKOUT0(soc_videooverlaysoc_hdmi_in0_mmcm_clk0_o),
	.CLKOUT2(soc_videooverlaysoc_hdmi_in0_mmcm_clk2_o),
	.DO(soc_videooverlaysoc_hdmi_in0_mmcm_dat_o_r_status),
	.DRDY(soc_videooverlaysoc_hdmi_in0_mmcm_drdy_o),
	.LOCKED(soc_videooverlaysoc_hdmi_in0_mmcm_locked_o)
);

BUFG BUFG_9(
	.I(soc_videooverlaysoc_hdmi_in0_mmcm_clk0_o),
	.O(pix_o_clk)
);

BUFG BUFG_10(
	.I(soc_videooverlaysoc_hdmi_in0_mmcm_clk2_o),
	.O(pix5x_o_clk)
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT(
	.I(hdmi_in0_data0_p),
	.IB(hdmi_in0_data0_n),
	.O(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_i_nodelay),
	.OB(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_32 (
	.C(hdmi_in0_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_master_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_master_inc),
	.LD(soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_32 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(hdmi_in0_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_i_delayed),
	.RST(hdmi_in0_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_33 (
	.C(hdmi_in0_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_slave_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_slave_inc),
	.LD(soc_videooverlaysoc_hdmi_in0_s7datacapture0_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_33 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(hdmi_in0_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_i_delayed),
	.RST(hdmi_in0_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in0_s7datacapture0_serdes_s_q[0])
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT_1(
	.I(hdmi_in0_data1_p),
	.IB(hdmi_in0_data1_n),
	.O(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_i_nodelay),
	.OB(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_34 (
	.C(hdmi_in0_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_master_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_master_inc),
	.LD(soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_34 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(hdmi_in0_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_i_delayed),
	.RST(hdmi_in0_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_35 (
	.C(hdmi_in0_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_slave_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_slave_inc),
	.LD(soc_videooverlaysoc_hdmi_in0_s7datacapture1_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_35 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(hdmi_in0_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_i_delayed),
	.RST(hdmi_in0_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in0_s7datacapture1_serdes_s_q[0])
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT_2(
	.I(hdmi_in0_data2_p),
	.IB(hdmi_in0_data2_n),
	.O(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_i_nodelay),
	.OB(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_36 (
	.C(hdmi_in0_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_master_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_master_inc),
	.LD(soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_36 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(hdmi_in0_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_i_delayed),
	.RST(hdmi_in0_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_37 (
	.C(hdmi_in0_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_slave_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_slave_inc),
	.LD(soc_videooverlaysoc_hdmi_in0_s7datacapture2_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_37 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(hdmi_in0_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_i_delayed),
	.RST(hdmi_in0_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in0_s7datacapture2_serdes_s_q[0])
);

reg [20:0] storage_10[0:7];
reg [2:0] memadr_6;
always @(posedge hdmi_in0_pix_clk) begin
	if (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_we)
		storage_10[soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_adr] <= soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_dat_w;
	memadr_6 <= soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_wrport_dat_r = storage_10[memadr_6];
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_rdport_dat_r = storage_10[soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer0_rdport_adr];

reg [20:0] storage_11[0:7];
reg [2:0] memadr_7;
always @(posedge hdmi_in0_pix_clk) begin
	if (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_we)
		storage_11[soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_adr] <= soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_dat_w;
	memadr_7 <= soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_wrport_dat_r = storage_11[memadr_7];
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_rdport_dat_r = storage_11[soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer1_rdport_adr];

reg [20:0] storage_12[0:7];
reg [2:0] memadr_8;
always @(posedge hdmi_in0_pix_clk) begin
	if (soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_we)
		storage_12[soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_adr] <= soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_dat_w;
	memadr_8 <= soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_wrport_dat_r = storage_12[memadr_8];
assign soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_rdport_dat_r = storage_12[soc_videooverlaysoc_hdmi_in0_chansync_syncbuffer2_rdport_adr];

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_65 (
	.CLK(pix5x_o_clk),
	.CLKDIV(pix_o_clk),
	.D1(soc_videooverlaysoc_hdmi_out0_clk_gen_data1[0]),
	.D2(soc_videooverlaysoc_hdmi_out0_clk_gen_data1[1]),
	.D3(soc_videooverlaysoc_hdmi_out0_clk_gen_data1[2]),
	.D4(soc_videooverlaysoc_hdmi_out0_clk_gen_data1[3]),
	.D5(soc_videooverlaysoc_hdmi_out0_clk_gen_data1[4]),
	.D6(soc_videooverlaysoc_hdmi_out0_clk_gen_data1[5]),
	.D7(soc_videooverlaysoc_hdmi_out0_clk_gen_data1[6]),
	.D8(soc_videooverlaysoc_hdmi_out0_clk_gen_data1[7]),
	.OCE(soc_videooverlaysoc_hdmi_out0_clk_gen_ce),
	.RST(pix_o_rst),
	.SHIFTIN1(soc_videooverlaysoc_hdmi_out0_clk_gen_shift[0]),
	.SHIFTIN2(soc_videooverlaysoc_hdmi_out0_clk_gen_shift[1]),
	.TCE(1'd0),
	.OQ(soc_videooverlaysoc_hdmi_out0_clk_gen_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_66 (
	.CLK(pix5x_o_clk),
	.CLKDIV(pix_o_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(soc_videooverlaysoc_hdmi_out0_clk_gen_data1[8]),
	.D4(soc_videooverlaysoc_hdmi_out0_clk_gen_data1[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(soc_videooverlaysoc_hdmi_out0_clk_gen_ce),
	.RST(pix_o_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(soc_videooverlaysoc_hdmi_out0_clk_gen_shift[0]),
	.SHIFTOUT2(soc_videooverlaysoc_hdmi_out0_clk_gen_shift[1])
);

OBUFDS OBUFDS_1(
	.I(soc_videooverlaysoc_hdmi_out0_clk_gen_pad_se),
	.O(hdmi_out0_clk_p),
	.OB(hdmi_out0_clk_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_67 (
	.CLK(pix5x_o_clk),
	.CLKDIV(pix_o_clk),
	.D1(soc_videooverlaysoc_hdmi_out0_phy_es0_data1[0]),
	.D2(soc_videooverlaysoc_hdmi_out0_phy_es0_data1[1]),
	.D3(soc_videooverlaysoc_hdmi_out0_phy_es0_data1[2]),
	.D4(soc_videooverlaysoc_hdmi_out0_phy_es0_data1[3]),
	.D5(soc_videooverlaysoc_hdmi_out0_phy_es0_data1[4]),
	.D6(soc_videooverlaysoc_hdmi_out0_phy_es0_data1[5]),
	.D7(soc_videooverlaysoc_hdmi_out0_phy_es0_data1[6]),
	.D8(soc_videooverlaysoc_hdmi_out0_phy_es0_data1[7]),
	.OCE(soc_videooverlaysoc_hdmi_out0_phy_es0_ce),
	.RST(pix_o_rst),
	.SHIFTIN1(soc_videooverlaysoc_hdmi_out0_phy_es0_shift[0]),
	.SHIFTIN2(soc_videooverlaysoc_hdmi_out0_phy_es0_shift[1]),
	.TCE(1'd0),
	.OQ(soc_videooverlaysoc_hdmi_out0_phy_es0_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_68 (
	.CLK(pix5x_o_clk),
	.CLKDIV(pix_o_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(soc_videooverlaysoc_hdmi_out0_phy_es0_data1[8]),
	.D4(soc_videooverlaysoc_hdmi_out0_phy_es0_data1[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(soc_videooverlaysoc_hdmi_out0_phy_es0_ce),
	.RST(pix_o_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(soc_videooverlaysoc_hdmi_out0_phy_es0_shift[0]),
	.SHIFTOUT2(soc_videooverlaysoc_hdmi_out0_phy_es0_shift[1])
);

OBUFDS OBUFDS_2(
	.I(soc_videooverlaysoc_hdmi_out0_phy_es0_pad_se),
	.O(hdmi_out0_data0_p),
	.OB(hdmi_out0_data0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_69 (
	.CLK(pix5x_o_clk),
	.CLKDIV(pix_o_clk),
	.D1(soc_videooverlaysoc_hdmi_out0_phy_es1_data1[0]),
	.D2(soc_videooverlaysoc_hdmi_out0_phy_es1_data1[1]),
	.D3(soc_videooverlaysoc_hdmi_out0_phy_es1_data1[2]),
	.D4(soc_videooverlaysoc_hdmi_out0_phy_es1_data1[3]),
	.D5(soc_videooverlaysoc_hdmi_out0_phy_es1_data1[4]),
	.D6(soc_videooverlaysoc_hdmi_out0_phy_es1_data1[5]),
	.D7(soc_videooverlaysoc_hdmi_out0_phy_es1_data1[6]),
	.D8(soc_videooverlaysoc_hdmi_out0_phy_es1_data1[7]),
	.OCE(soc_videooverlaysoc_hdmi_out0_phy_es1_ce),
	.RST(pix_o_rst),
	.SHIFTIN1(soc_videooverlaysoc_hdmi_out0_phy_es1_shift[0]),
	.SHIFTIN2(soc_videooverlaysoc_hdmi_out0_phy_es1_shift[1]),
	.TCE(1'd0),
	.OQ(soc_videooverlaysoc_hdmi_out0_phy_es1_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_70 (
	.CLK(pix5x_o_clk),
	.CLKDIV(pix_o_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(soc_videooverlaysoc_hdmi_out0_phy_es1_data1[8]),
	.D4(soc_videooverlaysoc_hdmi_out0_phy_es1_data1[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(soc_videooverlaysoc_hdmi_out0_phy_es1_ce),
	.RST(pix_o_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(soc_videooverlaysoc_hdmi_out0_phy_es1_shift[0]),
	.SHIFTOUT2(soc_videooverlaysoc_hdmi_out0_phy_es1_shift[1])
);

OBUFDS OBUFDS_3(
	.I(soc_videooverlaysoc_hdmi_out0_phy_es1_pad_se),
	.O(hdmi_out0_data1_p),
	.OB(hdmi_out0_data1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_71 (
	.CLK(pix5x_o_clk),
	.CLKDIV(pix_o_clk),
	.D1(soc_videooverlaysoc_hdmi_out0_phy_es2_data1[0]),
	.D2(soc_videooverlaysoc_hdmi_out0_phy_es2_data1[1]),
	.D3(soc_videooverlaysoc_hdmi_out0_phy_es2_data1[2]),
	.D4(soc_videooverlaysoc_hdmi_out0_phy_es2_data1[3]),
	.D5(soc_videooverlaysoc_hdmi_out0_phy_es2_data1[4]),
	.D6(soc_videooverlaysoc_hdmi_out0_phy_es2_data1[5]),
	.D7(soc_videooverlaysoc_hdmi_out0_phy_es2_data1[6]),
	.D8(soc_videooverlaysoc_hdmi_out0_phy_es2_data1[7]),
	.OCE(soc_videooverlaysoc_hdmi_out0_phy_es2_ce),
	.RST(pix_o_rst),
	.SHIFTIN1(soc_videooverlaysoc_hdmi_out0_phy_es2_shift[0]),
	.SHIFTIN2(soc_videooverlaysoc_hdmi_out0_phy_es2_shift[1]),
	.TCE(1'd0),
	.OQ(soc_videooverlaysoc_hdmi_out0_phy_es2_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_72 (
	.CLK(pix5x_o_clk),
	.CLKDIV(pix_o_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(soc_videooverlaysoc_hdmi_out0_phy_es2_data1[8]),
	.D4(soc_videooverlaysoc_hdmi_out0_phy_es2_data1[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(soc_videooverlaysoc_hdmi_out0_phy_es2_ce),
	.RST(pix_o_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(soc_videooverlaysoc_hdmi_out0_phy_es2_shift[0]),
	.SHIFTOUT2(soc_videooverlaysoc_hdmi_out0_phy_es2_shift[1])
);

OBUFDS OBUFDS_4(
	.I(soc_videooverlaysoc_hdmi_out0_phy_es2_pad_se),
	.O(hdmi_out0_data2_p),
	.OB(hdmi_out0_data2_n)
);

reg [7:0] edid_mem_1[0:255];
reg [7:0] memadr_9;
reg [7:0] memadr_10;
always @(posedge sys_clk) begin
	memadr_9 <= soc_videooverlaysoc_hdmi_in1_edid_adr;
end

always @(posedge sys_clk) begin
	if (vns_videooverlaysoc_sram1_we)
		edid_mem_1[vns_videooverlaysoc_sram1_adr] <= vns_videooverlaysoc_sram1_dat_w;
	memadr_10 <= vns_videooverlaysoc_sram1_adr;
end

assign soc_videooverlaysoc_hdmi_in1_edid_dat_r = edid_mem_1[memadr_9];
assign vns_videooverlaysoc_sram1_dat_r = edid_mem_1[memadr_10];

initial begin
	$readmemh("edid_mem_1.init", edid_mem_1);
end

assign hdmi_in1_sda = soc_videooverlaysoc_hdmi_in1_edid_sda_drv_reg ? 1'd0 : 1'bz;
assign soc_videooverlaysoc_hdmi_in1_edid_sda_i_async = hdmi_in1_sda;

IBUFDS_DIFF_OUT hdmi_in_ibufds_1(
	.I(hdmi_in1_clk_p),
	.IB(hdmi_in1_clk_n),
	.O(soc_videooverlaysoc_hdmi_in1_clk_input)
);

BUFR BUFR_1(
	.I(soc_videooverlaysoc_hdmi_in1_clk_input),
	.O(soc_videooverlaysoc_hdmi_in1_clk_input_bufr)
);

MMCME2_ADV #(
	.BANDWIDTH("OPTIMIZED"),
	.CLKFBOUT_MULT_F(5.0),
	.CLKFBOUT_PHASE(0.0),
	.CLKIN1_PERIOD(6.734),
	.CLKOUT0_DIVIDE_F(3'd5),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(3'd4),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(1'd1),
	.CLKOUT2_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01)
) MMCME2_ADV_1 (
	.CLKFBIN(soc_videooverlaysoc_hdmi_in1_mmcm_fb_o),
	.CLKIN1(soc_videooverlaysoc_hdmi_in1_clk_input_bufr),
	.DADDR(soc_videooverlaysoc_hdmi_in1_mmcm_adr_storage),
	.DCLK(sys_clk),
	.DEN((soc_videooverlaysoc_hdmi_in1_mmcm_read_re | soc_videooverlaysoc_hdmi_in1_mmcm_write_re)),
	.DI(soc_videooverlaysoc_hdmi_in1_mmcm_dat_w_storage),
	.DWE(soc_videooverlaysoc_hdmi_in1_mmcm_write_re),
	.RST(soc_videooverlaysoc_hdmi_in1_mmcm_reset_storage),
	.CLKFBOUT(soc_videooverlaysoc_hdmi_in1_mmcm_fb),
	.CLKOUT0(soc_videooverlaysoc_hdmi_in1_mmcm_clk0),
	.CLKOUT1(soc_videooverlaysoc_hdmi_in1_mmcm_clk1),
	.CLKOUT2(soc_videooverlaysoc_hdmi_in1_mmcm_clk2),
	.DO(soc_videooverlaysoc_hdmi_in1_mmcm_dat_r_status),
	.DRDY(soc_videooverlaysoc_hdmi_in1_mmcm_drdy),
	.LOCKED(soc_videooverlaysoc_hdmi_in1_mmcm_locked)
);

BUFG BUFG_11(
	.I(soc_videooverlaysoc_hdmi_in1_mmcm_clk0),
	.O(hdmi_in1_pix_clk)
);

BUFG BUFG_12(
	.I(soc_videooverlaysoc_hdmi_in1_mmcm_clk1),
	.O(hdmi_in1_pix1p25x_clk)
);

BUFIO BUFIO_1(
	.I(soc_videooverlaysoc_hdmi_in1_mmcm_clk2),
	.O(hdmi_in1_pix5x_clk)
);

BUFG BUFG_13(
	.I(soc_videooverlaysoc_hdmi_in1_mmcm_fb),
	.O(soc_videooverlaysoc_hdmi_in1_mmcm_fb_o)
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT_3(
	.I(hdmi_in1_data0_p),
	.IB(hdmi_in1_data0_n),
	.O(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_i_nodelay),
	.OB(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_38 (
	.C(hdmi_in1_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_master_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_master_inc),
	.LD(soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_38 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in1_pix5x_clk),
	.CLKB((~hdmi_in1_pix5x_clk)),
	.CLKDIV(hdmi_in1_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_i_delayed),
	.RST(hdmi_in1_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_39 (
	.C(hdmi_in1_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_slave_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_slave_inc),
	.LD(soc_videooverlaysoc_hdmi_in1_s7datacapture0_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_39 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in1_pix5x_clk),
	.CLKB((~hdmi_in1_pix5x_clk)),
	.CLKDIV(hdmi_in1_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_i_delayed),
	.RST(hdmi_in1_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in1_s7datacapture0_serdes_s_q[0])
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT_4(
	.I(hdmi_in1_data1_p),
	.IB(hdmi_in1_data1_n),
	.O(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_i_nodelay),
	.OB(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_40 (
	.C(hdmi_in1_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_master_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_master_inc),
	.LD(soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_40 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in1_pix5x_clk),
	.CLKB((~hdmi_in1_pix5x_clk)),
	.CLKDIV(hdmi_in1_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_i_delayed),
	.RST(hdmi_in1_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_41 (
	.C(hdmi_in1_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_slave_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_slave_inc),
	.LD(soc_videooverlaysoc_hdmi_in1_s7datacapture1_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_41 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in1_pix5x_clk),
	.CLKB((~hdmi_in1_pix5x_clk)),
	.CLKDIV(hdmi_in1_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_i_delayed),
	.RST(hdmi_in1_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in1_s7datacapture1_serdes_s_q[0])
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT_5(
	.I(hdmi_in1_data2_p),
	.IB(hdmi_in1_data2_n),
	.O(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_i_nodelay),
	.OB(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_42 (
	.C(hdmi_in1_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_master_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_master_inc),
	.LD(soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_42 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in1_pix5x_clk),
	.CLKB((~hdmi_in1_pix5x_clk)),
	.CLKDIV(hdmi_in1_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_i_delayed),
	.RST(hdmi_in1_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_43 (
	.C(hdmi_in1_pix1p25x_clk),
	.CE(soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_slave_ce),
	.IDATAIN(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_i_nodelay),
	.INC(soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_slave_inc),
	.LD(soc_videooverlaysoc_hdmi_in1_s7datacapture2_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_43 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in1_pix5x_clk),
	.CLKB((~hdmi_in1_pix5x_clk)),
	.CLKDIV(hdmi_in1_pix1p25x_clk),
	.DDLY(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_i_delayed),
	.RST(hdmi_in1_pix1p25x_rst),
	.Q1(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_q[7]),
	.Q2(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_q[6]),
	.Q3(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_q[5]),
	.Q4(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_q[4]),
	.Q5(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_q[3]),
	.Q6(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_q[2]),
	.Q7(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_q[1]),
	.Q8(soc_videooverlaysoc_hdmi_in1_s7datacapture2_serdes_s_q[0])
);

reg [20:0] storage_13[0:7];
reg [2:0] memadr_11;
always @(posedge hdmi_in1_pix_clk) begin
	if (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_we)
		storage_13[soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_adr] <= soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_dat_w;
	memadr_11 <= soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_adr;
end

always @(posedge hdmi_in1_pix_clk) begin
end

assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_wrport_dat_r = storage_13[memadr_11];
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_rdport_dat_r = storage_13[soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer0_rdport_adr];

reg [20:0] storage_14[0:7];
reg [2:0] memadr_12;
always @(posedge hdmi_in1_pix_clk) begin
	if (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_we)
		storage_14[soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_adr] <= soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_dat_w;
	memadr_12 <= soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_adr;
end

always @(posedge hdmi_in1_pix_clk) begin
end

assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_wrport_dat_r = storage_14[memadr_12];
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_rdport_dat_r = storage_14[soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer1_rdport_adr];

reg [20:0] storage_15[0:7];
reg [2:0] memadr_13;
always @(posedge hdmi_in1_pix_clk) begin
	if (soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_we)
		storage_15[soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_adr] <= soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_dat_w;
	memadr_13 <= soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_adr;
end

always @(posedge hdmi_in1_pix_clk) begin
end

assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_wrport_dat_r = storage_15[memadr_13];
assign soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_rdport_dat_r = storage_15[soc_videooverlaysoc_hdmi_in1_chansync_syncbuffer2_rdport_adr];

reg [258:0] storage_16[0:1023];
reg [9:0] memadr_14;
reg [9:0] memadr_15;
always @(posedge hdmi_in1_pix_clk) begin
	if (soc_videooverlaysoc_hdmi_in1_frame_wrport_we)
		storage_16[soc_videooverlaysoc_hdmi_in1_frame_wrport_adr] <= soc_videooverlaysoc_hdmi_in1_frame_wrport_dat_w;
	memadr_14 <= soc_videooverlaysoc_hdmi_in1_frame_wrport_adr;
end

always @(posedge sys_clk) begin
	memadr_15 <= soc_videooverlaysoc_hdmi_in1_frame_rdport_adr;
end

assign soc_videooverlaysoc_hdmi_in1_frame_wrport_dat_r = storage_16[memadr_14];
assign soc_videooverlaysoc_hdmi_in1_frame_rdport_dat_r = storage_16[memadr_15];

reg [257:0] storage_17[0:15];
reg [257:0] memdat_12;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_we)
		storage_17[soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_adr] <= soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_dat_w;
	memdat_12 <= storage_17[soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign soc_videooverlaysoc_hdmi_in1_dma_fifo_wrport_dat_r = memdat_12;
assign soc_videooverlaysoc_hdmi_in1_dma_fifo_rdport_dat_r = storage_17[soc_videooverlaysoc_hdmi_in1_dma_fifo_rdport_adr];

reg [26:0] storage_18[0:3];
reg [1:0] memadr_16;
reg [1:0] memadr_17;
always @(posedge pix_o_clk) begin
	if (soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_we)
		storage_18[soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_adr] <= soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_dat_w;
	memadr_16 <= soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
	memadr_17 <= soc_videooverlaysoc_out_dram_port_cmd_fifo_rdport_adr;
end

assign soc_videooverlaysoc_out_dram_port_cmd_fifo_wrport_dat_r = storage_18[memadr_16];
assign soc_videooverlaysoc_out_dram_port_cmd_fifo_rdport_dat_r = storage_18[memadr_17];

reg [257:0] storage_19[0:15];
reg [3:0] memadr_18;
reg [3:0] memadr_19;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_we)
		storage_19[soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_adr] <= soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_dat_w;
	memadr_18 <= soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_adr;
end

always @(posedge pix_o_clk) begin
	memadr_19 <= soc_videooverlaysoc_out_dram_port_rdata_fifo_rdport_adr;
end

assign soc_videooverlaysoc_out_dram_port_rdata_fifo_wrport_dat_r = storage_19[memadr_18];
assign soc_videooverlaysoc_out_dram_port_rdata_fifo_rdport_dat_r = storage_19[memadr_19];

reg [9:0] storage_20[0:3];
reg [9:0] memdat_13;
always @(posedge pix_o_clk) begin
	if (soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_we)
		storage_20[soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_adr] <= soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_dat_w;
	memdat_13 <= storage_20[soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_adr];
end

always @(posedge pix_o_clk) begin
end

assign soc_videooverlaysoc_out_dram_port_cmd_buffer_wrport_dat_r = memdat_13;
assign soc_videooverlaysoc_out_dram_port_cmd_buffer_rdport_dat_r = storage_20[soc_videooverlaysoc_out_dram_port_cmd_buffer_rdport_adr];

reg [161:0] storage_21[0:1];
reg [0:0] memadr_20;
reg [0:0] memadr_21;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_we)
		storage_21[soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_adr] <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_dat_w;
	memadr_20 <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_adr;
end

always @(posedge pix_o_clk) begin
	memadr_21 <= soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_rdport_adr;
end

assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_wrport_dat_r = storage_21[memadr_20];
assign soc_videooverlaysoc_hdmi_core_out0_initiator_cdc_rdport_dat_r = storage_21[memadr_21];

reg [33:0] storage_22[0:1023];
reg [33:0] memdat_14;
reg [33:0] memdat_15;
always @(posedge pix_o_clk) begin
	if (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_we)
		storage_22[soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_adr] <= soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_dat_w;
	memdat_14 <= storage_22[soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_adr];
end

always @(posedge pix_o_clk) begin
	if (soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_rdport_re)
		memdat_15 <= storage_22[soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_rdport_adr];
end

assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_wrport_dat_r = memdat_14;
assign soc_videooverlaysoc_hdmi_core_out0_dmareader_fifo_rdport_dat_r = memdat_15;

i2c_snoop i2c_snoop(
	.SCL((~hdmi_in0_scl)),
	.SDA((~hdmi_in0_sda)),
	.clk(eth_clk),
	.i2c_snoop_addr(7'd116),
	.reg_addr(soc_videooverlaysoc_i2c_snoop_storage),
	.reset(eth_rst),
	.Aksv14_write(soc_videooverlaysoc_i2c_snoop_Aksv14_write),
	.An(soc_videooverlaysoc_i2c_snoop_An),
	.reg_dout(soc_videooverlaysoc_i2c_snoop_reg_dout)
);

hdcp_mod hdcp_mod(
	.Aksv14_write(soc_videooverlaysoc_hdcp_Aksv14_write),
	.An(soc_videooverlaysoc_hdcp_An),
	.Km(soc_videooverlaysoc_hdcp_Km_storage),
	.Km_valid(soc_videooverlaysoc_hdcp_Km_valid_storage),
	.clk(pix_o_clk),
	.ctl_code(soc_videooverlaysoc_hdcp_ctl_code),
	.de(soc_videooverlaysoc_hdmi_in0_timing_payload_de),
	.hdcp_ena(soc_videooverlaysoc_hdcp_hdcp_ena),
	.hpd(soc_videooverlaysoc_hdcp_hpd),
	.hsync(soc_videooverlaysoc_hdmi_in0_timing_payload_hsync),
	.line_end(soc_videooverlaysoc_hdcp_line_end),
	.rst(pix_o_rst),
	.vsync(soc_videooverlaysoc_hdmi_in0_timing_payload_vsync),
	.cipher_stream(soc_videooverlaysoc_hdcp_cipher_stream),
	.stream_ready(soc_videooverlaysoc_hdcp_stream_ready)
);

assign rmii_eth_mdio = soc_videooverlaysoc_phy_data_oe ? soc_videooverlaysoc_phy_data_w : 1'bz;
assign soc_videooverlaysoc_phy_data_r = rmii_eth_mdio;

reg [11:0] storage_23[0:4];
reg [11:0] memdat_16;
always @(posedge eth_rx_clk) begin
	if (soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_we)
		storage_23[soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_adr] <= soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_dat_w;
	memdat_16 <= storage_23[soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_adr];
end

always @(posedge eth_rx_clk) begin
end

assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_wrport_dat_r = memdat_16;
assign soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_rdport_dat_r = storage_23[soc_videooverlaysoc_core_mac_crc32_checker_syncfifo_rdport_adr];

reg [11:0] storage_24[0:63];
reg [5:0] memadr_22;
reg [5:0] memadr_23;
always @(posedge eth_clk) begin
	if (soc_videooverlaysoc_core_mac_tx_cdc_wrport_we)
		storage_24[soc_videooverlaysoc_core_mac_tx_cdc_wrport_adr] <= soc_videooverlaysoc_core_mac_tx_cdc_wrport_dat_w;
	memadr_22 <= soc_videooverlaysoc_core_mac_tx_cdc_wrport_adr;
end

always @(posedge eth_tx_clk) begin
	memadr_23 <= soc_videooverlaysoc_core_mac_tx_cdc_rdport_adr;
end

assign soc_videooverlaysoc_core_mac_tx_cdc_wrport_dat_r = storage_24[memadr_22];
assign soc_videooverlaysoc_core_mac_tx_cdc_rdport_dat_r = storage_24[memadr_23];

reg [11:0] storage_25[0:63];
reg [5:0] memadr_24;
reg [5:0] memadr_25;
always @(posedge eth_rx_clk) begin
	if (soc_videooverlaysoc_core_mac_rx_cdc_wrport_we)
		storage_25[soc_videooverlaysoc_core_mac_rx_cdc_wrport_adr] <= soc_videooverlaysoc_core_mac_rx_cdc_wrport_dat_w;
	memadr_24 <= soc_videooverlaysoc_core_mac_rx_cdc_wrport_adr;
end

always @(posedge eth_clk) begin
	memadr_25 <= soc_videooverlaysoc_core_mac_rx_cdc_rdport_adr;
end

assign soc_videooverlaysoc_core_mac_rx_cdc_wrport_dat_r = storage_25[memadr_24];
assign soc_videooverlaysoc_core_mac_rx_cdc_rdport_dat_r = storage_25[memadr_25];

reg [122:0] storage_26[0:127];
reg [122:0] memdat_17;
reg [122:0] memdat_18;
always @(posedge eth_clk) begin
	if (soc_videooverlaysoc_core_icmp_echo_buffer_wrport_we)
		storage_26[soc_videooverlaysoc_core_icmp_echo_buffer_wrport_adr] <= soc_videooverlaysoc_core_icmp_echo_buffer_wrport_dat_w;
	memdat_17 <= storage_26[soc_videooverlaysoc_core_icmp_echo_buffer_wrport_adr];
end

always @(posedge eth_clk) begin
	if (soc_videooverlaysoc_core_icmp_echo_buffer_rdport_re)
		memdat_18 <= storage_26[soc_videooverlaysoc_core_icmp_echo_buffer_rdport_adr];
end

assign soc_videooverlaysoc_core_icmp_echo_buffer_wrport_dat_r = memdat_17;
assign soc_videooverlaysoc_core_icmp_echo_buffer_rdport_dat_r = memdat_18;

reg [117:0] storage_27[0:3];
reg [1:0] memadr_26;
reg [1:0] memadr_27;
always @(posedge etherbone_clk) begin
	if (soc_videooverlaysoc_packet_tx_cdc_wrport_we)
		storage_27[soc_videooverlaysoc_packet_tx_cdc_wrport_adr] <= soc_videooverlaysoc_packet_tx_cdc_wrport_dat_w;
	memadr_26 <= soc_videooverlaysoc_packet_tx_cdc_wrport_adr;
end

always @(posedge eth_clk) begin
	memadr_27 <= soc_videooverlaysoc_packet_tx_cdc_rdport_adr;
end

assign soc_videooverlaysoc_packet_tx_cdc_wrport_dat_r = storage_27[memadr_26];
assign soc_videooverlaysoc_packet_tx_cdc_rdport_dat_r = storage_27[memadr_27];

reg [117:0] storage_28[0:3];
reg [1:0] memadr_28;
reg [1:0] memadr_29;
always @(posedge eth_clk) begin
	if (soc_videooverlaysoc_packet_rx_cdc_wrport_we)
		storage_28[soc_videooverlaysoc_packet_rx_cdc_wrport_adr] <= soc_videooverlaysoc_packet_rx_cdc_wrport_dat_w;
	memadr_28 <= soc_videooverlaysoc_packet_rx_cdc_wrport_adr;
end

always @(posedge etherbone_clk) begin
	memadr_29 <= soc_videooverlaysoc_packet_rx_cdc_rdport_adr;
end

assign soc_videooverlaysoc_packet_rx_cdc_wrport_dat_r = storage_28[memadr_28];
assign soc_videooverlaysoc_packet_rx_cdc_rdport_dat_r = storage_28[memadr_29];

reg [67:0] storage_29[0:3];
reg [67:0] memdat_19;
reg [67:0] memdat_20;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_record_receiver_fifo_wrport_we)
		storage_29[soc_videooverlaysoc_record_receiver_fifo_wrport_adr] <= soc_videooverlaysoc_record_receiver_fifo_wrport_dat_w;
	memdat_19 <= storage_29[soc_videooverlaysoc_record_receiver_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_record_receiver_fifo_rdport_re)
		memdat_20 <= storage_29[soc_videooverlaysoc_record_receiver_fifo_rdport_adr];
end

assign soc_videooverlaysoc_record_receiver_fifo_wrport_dat_r = memdat_19;
assign soc_videooverlaysoc_record_receiver_fifo_rdport_dat_r = memdat_20;

reg [110:0] storage_30[0:3];
reg [110:0] memdat_21;
reg [110:0] memdat_22;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_record_sender_fifo_wrport_we)
		storage_30[soc_videooverlaysoc_record_sender_fifo_wrport_adr] <= soc_videooverlaysoc_record_sender_fifo_wrport_dat_w;
	memdat_21 <= storage_30[soc_videooverlaysoc_record_sender_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_record_sender_fifo_rdport_re)
		memdat_22 <= storage_30[soc_videooverlaysoc_record_sender_fifo_rdport_adr];
end

assign soc_videooverlaysoc_record_sender_fifo_wrport_dat_r = memdat_21;
assign soc_videooverlaysoc_record_sender_fifo_rdport_dat_r = memdat_22;

reg [7:0] data_mem_grain0[0:255];
reg [7:0] memadr_30;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[0])
		data_mem_grain0[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[7:0];
	memadr_30 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[7:0] = data_mem_grain0[memadr_30];

reg [7:0] data_mem_grain1[0:255];
reg [7:0] memadr_31;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[1])
		data_mem_grain1[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[15:8];
	memadr_31 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[15:8] = data_mem_grain1[memadr_31];

reg [7:0] data_mem_grain2[0:255];
reg [7:0] memadr_32;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[2])
		data_mem_grain2[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[23:16];
	memadr_32 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[23:16] = data_mem_grain2[memadr_32];

reg [7:0] data_mem_grain3[0:255];
reg [7:0] memadr_33;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[3])
		data_mem_grain3[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[31:24];
	memadr_33 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[31:24] = data_mem_grain3[memadr_33];

reg [7:0] data_mem_grain4[0:255];
reg [7:0] memadr_34;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[4])
		data_mem_grain4[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[39:32];
	memadr_34 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[39:32] = data_mem_grain4[memadr_34];

reg [7:0] data_mem_grain5[0:255];
reg [7:0] memadr_35;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[5])
		data_mem_grain5[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[47:40];
	memadr_35 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[47:40] = data_mem_grain5[memadr_35];

reg [7:0] data_mem_grain6[0:255];
reg [7:0] memadr_36;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[6])
		data_mem_grain6[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[55:48];
	memadr_36 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[55:48] = data_mem_grain6[memadr_36];

reg [7:0] data_mem_grain7[0:255];
reg [7:0] memadr_37;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[7])
		data_mem_grain7[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[63:56];
	memadr_37 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[63:56] = data_mem_grain7[memadr_37];

reg [7:0] data_mem_grain8[0:255];
reg [7:0] memadr_38;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[8])
		data_mem_grain8[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[71:64];
	memadr_38 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[71:64] = data_mem_grain8[memadr_38];

reg [7:0] data_mem_grain9[0:255];
reg [7:0] memadr_39;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[9])
		data_mem_grain9[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[79:72];
	memadr_39 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[79:72] = data_mem_grain9[memadr_39];

reg [7:0] data_mem_grain10[0:255];
reg [7:0] memadr_40;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[10])
		data_mem_grain10[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[87:80];
	memadr_40 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[87:80] = data_mem_grain10[memadr_40];

reg [7:0] data_mem_grain11[0:255];
reg [7:0] memadr_41;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[11])
		data_mem_grain11[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[95:88];
	memadr_41 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[95:88] = data_mem_grain11[memadr_41];

reg [7:0] data_mem_grain12[0:255];
reg [7:0] memadr_42;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[12])
		data_mem_grain12[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[103:96];
	memadr_42 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[103:96] = data_mem_grain12[memadr_42];

reg [7:0] data_mem_grain13[0:255];
reg [7:0] memadr_43;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[13])
		data_mem_grain13[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[111:104];
	memadr_43 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[111:104] = data_mem_grain13[memadr_43];

reg [7:0] data_mem_grain14[0:255];
reg [7:0] memadr_44;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[14])
		data_mem_grain14[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[119:112];
	memadr_44 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[119:112] = data_mem_grain14[memadr_44];

reg [7:0] data_mem_grain15[0:255];
reg [7:0] memadr_45;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[15])
		data_mem_grain15[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[127:120];
	memadr_45 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[127:120] = data_mem_grain15[memadr_45];

reg [7:0] data_mem_grain16[0:255];
reg [7:0] memadr_46;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[16])
		data_mem_grain16[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[135:128];
	memadr_46 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[135:128] = data_mem_grain16[memadr_46];

reg [7:0] data_mem_grain17[0:255];
reg [7:0] memadr_47;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[17])
		data_mem_grain17[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[143:136];
	memadr_47 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[143:136] = data_mem_grain17[memadr_47];

reg [7:0] data_mem_grain18[0:255];
reg [7:0] memadr_48;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[18])
		data_mem_grain18[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[151:144];
	memadr_48 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[151:144] = data_mem_grain18[memadr_48];

reg [7:0] data_mem_grain19[0:255];
reg [7:0] memadr_49;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[19])
		data_mem_grain19[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[159:152];
	memadr_49 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[159:152] = data_mem_grain19[memadr_49];

reg [7:0] data_mem_grain20[0:255];
reg [7:0] memadr_50;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[20])
		data_mem_grain20[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[167:160];
	memadr_50 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[167:160] = data_mem_grain20[memadr_50];

reg [7:0] data_mem_grain21[0:255];
reg [7:0] memadr_51;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[21])
		data_mem_grain21[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[175:168];
	memadr_51 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[175:168] = data_mem_grain21[memadr_51];

reg [7:0] data_mem_grain22[0:255];
reg [7:0] memadr_52;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[22])
		data_mem_grain22[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[183:176];
	memadr_52 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[183:176] = data_mem_grain22[memadr_52];

reg [7:0] data_mem_grain23[0:255];
reg [7:0] memadr_53;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[23])
		data_mem_grain23[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[191:184];
	memadr_53 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[191:184] = data_mem_grain23[memadr_53];

reg [7:0] data_mem_grain24[0:255];
reg [7:0] memadr_54;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[24])
		data_mem_grain24[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[199:192];
	memadr_54 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[199:192] = data_mem_grain24[memadr_54];

reg [7:0] data_mem_grain25[0:255];
reg [7:0] memadr_55;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[25])
		data_mem_grain25[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[207:200];
	memadr_55 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[207:200] = data_mem_grain25[memadr_55];

reg [7:0] data_mem_grain26[0:255];
reg [7:0] memadr_56;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[26])
		data_mem_grain26[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[215:208];
	memadr_56 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[215:208] = data_mem_grain26[memadr_56];

reg [7:0] data_mem_grain27[0:255];
reg [7:0] memadr_57;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[27])
		data_mem_grain27[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[223:216];
	memadr_57 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[223:216] = data_mem_grain27[memadr_57];

reg [7:0] data_mem_grain28[0:255];
reg [7:0] memadr_58;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[28])
		data_mem_grain28[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[231:224];
	memadr_58 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[231:224] = data_mem_grain28[memadr_58];

reg [7:0] data_mem_grain29[0:255];
reg [7:0] memadr_59;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[29])
		data_mem_grain29[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[239:232];
	memadr_59 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[239:232] = data_mem_grain29[memadr_59];

reg [7:0] data_mem_grain30[0:255];
reg [7:0] memadr_60;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[30])
		data_mem_grain30[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[247:240];
	memadr_60 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[247:240] = data_mem_grain30[memadr_60];

reg [7:0] data_mem_grain31[0:255];
reg [7:0] memadr_61;
always @(posedge sys_clk) begin
	if (soc_videooverlaysoc_videooverlaysoc_data_port_we[31])
		data_mem_grain31[soc_videooverlaysoc_videooverlaysoc_data_port_adr] <= soc_videooverlaysoc_videooverlaysoc_data_port_dat_w[255:248];
	memadr_61 <= soc_videooverlaysoc_videooverlaysoc_data_port_adr;
end

assign soc_videooverlaysoc_videooverlaysoc_data_port_dat_r[255:248] = data_mem_grain31[memadr_61];

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE (
	.C(sys_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl0),
	.Q(vns_xilinxasyncresetsynchronizerimpl0_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_1 (
	.C(sys_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl0_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl0),
	.Q(sys_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_2 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl1),
	.Q(vns_xilinxasyncresetsynchronizerimpl1_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_3 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl1_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl1),
	.Q(clk200_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_4 (
	.C(eth_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl2),
	.Q(vns_xilinxasyncresetsynchronizerimpl2_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_5 (
	.C(eth_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl2_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl2),
	.Q(eth_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_6 (
	.C(hdmi_in0_pix_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl3),
	.Q(vns_xilinxasyncresetsynchronizerimpl3_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_7 (
	.C(hdmi_in0_pix_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl3_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl3),
	.Q(hdmi_in0_pix_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_8 (
	.C(hdmi_in0_pix1p25x_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl4),
	.Q(vns_xilinxasyncresetsynchronizerimpl4_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_9 (
	.C(hdmi_in0_pix1p25x_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl4_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl4),
	.Q(hdmi_in0_pix1p25x_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_10 (
	.C(pix_o_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl5),
	.Q(vns_xilinxasyncresetsynchronizerimpl5_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_11 (
	.C(pix_o_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl5_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl5),
	.Q(pix_o_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_12 (
	.C(hdmi_in1_pix_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl6),
	.Q(vns_xilinxasyncresetsynchronizerimpl6_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_13 (
	.C(hdmi_in1_pix_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl6_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl6),
	.Q(hdmi_in1_pix_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_14 (
	.C(hdmi_in1_pix1p25x_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl7),
	.Q(vns_xilinxasyncresetsynchronizerimpl7_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_15 (
	.C(hdmi_in1_pix1p25x_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl7_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl7),
	.Q(hdmi_in1_pix1p25x_rst)
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(1'd0),
	.D2(1'd1),
	.R(1'd0),
	.S(1'd0),
	.Q(rmii_eth_clocks_ref_clk)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_16 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(soc_videooverlaysoc_phy_reset0),
	.Q(vns_xilinxasyncresetsynchronizerimpl8_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_17 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl8_rst_meta),
	.PRE(soc_videooverlaysoc_phy_reset0),
	.Q(eth_tx_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_18 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(soc_videooverlaysoc_phy_reset0),
	.Q(vns_xilinxasyncresetsynchronizerimpl9_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_19 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl9_rst_meta),
	.PRE(soc_videooverlaysoc_phy_reset0),
	.Q(eth_rx_rst)
);

endmodule
