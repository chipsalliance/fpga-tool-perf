// Copyright lowRISC contributors.
// Copyright 2018 ETH Zurich and University of Bologna, see also CREDITS.md.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

module ibex_prefetch_buffer (
	clk_i,
	rst_ni,
	req_i,
	branch_i,
	addr_i,
	ready_i,
	valid_o,
	rdata_o,
	addr_o,
	err_o,
	instr_req_o,
	instr_gnt_i,
	instr_addr_o,
	instr_rdata_i,
	instr_err_i,
	instr_pmp_err_i,
	instr_rvalid_i,
	busy_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire req_i;
	input wire branch_i;
	input wire [31:0] addr_i;
	input wire ready_i;
	output wire valid_o;
	output wire [31:0] rdata_o;
	output wire [31:0] addr_o;
	output wire err_o;
	output wire instr_req_o;
	input wire instr_gnt_i;
	output wire [31:0] instr_addr_o;
	input wire [31:0] instr_rdata_i;
	input wire instr_err_i;
	input wire instr_pmp_err_i;
	input wire instr_rvalid_i;
	output wire busy_o;
	localparam [31:0] NUM_REQS = 2;
	wire valid_new_req;
	wire valid_req;
	wire valid_req_d;
	reg valid_req_q;
	wire discard_req_d;
	reg discard_req_q;
	wire gnt_or_pmp_err;
	wire rvalid_or_pmp_err;
	wire [(NUM_REQS - 1):0] rdata_outstanding_n;
	wire [(NUM_REQS - 1):0] rdata_outstanding_s;
	reg [(NUM_REQS - 1):0] rdata_outstanding_q;
	wire [(NUM_REQS - 1):0] branch_discard_n;
	wire [(NUM_REQS - 1):0] branch_discard_s;
	reg [(NUM_REQS - 1):0] branch_discard_q;
	wire [(NUM_REQS - 1):0] rdata_pmp_err_n;
	wire [(NUM_REQS - 1):0] rdata_pmp_err_s;
	reg [(NUM_REQS - 1):0] rdata_pmp_err_q;
	wire [31:0] stored_addr_d;
	reg [31:0] stored_addr_q;
	wire stored_addr_en;
	wire [31:0] fetch_addr_d;
	reg [31:0] fetch_addr_q;
	wire fetch_addr_en;
	wire [31:0] instr_addr;
	wire [31:0] instr_addr_w_aligned;
	wire instr_or_pmp_err;
	wire fifo_valid;
	wire fifo_ready;
	wire fifo_clear;
	assign busy_o = (|rdata_outstanding_q | instr_req_o);
	assign instr_or_pmp_err = (instr_err_i | rdata_pmp_err_q[0]);
	assign fifo_clear = branch_i;
	ibex_fetch_fifo #(.NUM_REQS(NUM_REQS)) fifo_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clear_i(fifo_clear),
		.in_valid_i(fifo_valid),
		.in_addr_i(addr_i),
		.in_rdata_i(instr_rdata_i),
		.in_err_i(instr_or_pmp_err),
		.in_ready_o(fifo_ready),
		.out_valid_o(valid_o),
		.out_ready_i(ready_i),
		.out_rdata_o(rdata_o),
		.out_addr_o(addr_o),
		.out_err_o(err_o)
	);
	assign valid_new_req = ((req_i & (fifo_ready | branch_i)) & ~rdata_outstanding_q[(NUM_REQS - 1)]);
	assign valid_req = (valid_req_q | valid_new_req);
	assign gnt_or_pmp_err = (instr_gnt_i | instr_pmp_err_i);
	assign rvalid_or_pmp_err = (rdata_outstanding_q[0] & (instr_rvalid_i | rdata_pmp_err_q[0]));
	assign valid_req_d = (valid_req & ~gnt_or_pmp_err);
	assign discard_req_d = (valid_req_q & (branch_i | discard_req_q));
	assign stored_addr_en = ((valid_new_req & ~valid_req_q) & ~gnt_or_pmp_err);
	assign stored_addr_d = instr_addr;
	always @(posedge clk_i)
		if (stored_addr_en)
			stored_addr_q <= stored_addr_d;
	assign fetch_addr_en = (branch_i | (valid_new_req & ~valid_req_q));
	assign fetch_addr_d = ((branch_i ? addr_i : {fetch_addr_q[31:2], 2'b00}) + {{29 {1'b0}}, (valid_new_req & ~valid_req_q), 2'b00});
	always @(posedge clk_i)
		if (fetch_addr_en)
			fetch_addr_q <= fetch_addr_d;
	assign instr_addr = (valid_req_q ? stored_addr_q : (branch_i ? addr_i : fetch_addr_q));
	assign instr_addr_w_aligned = {instr_addr[31:2], 2'b00};
	generate
		genvar g_outstanding_reqs_i;
		for (g_outstanding_reqs_i = 0; (g_outstanding_reqs_i < NUM_REQS); g_outstanding_reqs_i = (g_outstanding_reqs_i + 1)) begin : g_outstanding_reqs
			if ((g_outstanding_reqs_i == 0)) begin : g_req0
				assign rdata_outstanding_n[g_outstanding_reqs_i] = ((valid_req & gnt_or_pmp_err) | rdata_outstanding_q[g_outstanding_reqs_i]);
				assign branch_discard_n[g_outstanding_reqs_i] = ((((valid_req & gnt_or_pmp_err) & discard_req_d) | (branch_i & rdata_outstanding_q[g_outstanding_reqs_i])) | branch_discard_q[g_outstanding_reqs_i]);
				assign rdata_pmp_err_n[g_outstanding_reqs_i] = (((valid_req & ~rdata_outstanding_q[g_outstanding_reqs_i]) & instr_pmp_err_i) | rdata_pmp_err_q[g_outstanding_reqs_i]);
			end
			else begin : g_reqtop
				assign rdata_outstanding_n[g_outstanding_reqs_i] = (((valid_req & gnt_or_pmp_err) & rdata_outstanding_q[(g_outstanding_reqs_i - 1)]) | rdata_outstanding_q[g_outstanding_reqs_i]);
				assign branch_discard_n[g_outstanding_reqs_i] = (((((valid_req & gnt_or_pmp_err) & discard_req_d) & rdata_outstanding_q[(g_outstanding_reqs_i - 1)]) | (branch_i & rdata_outstanding_q[g_outstanding_reqs_i])) | branch_discard_q[g_outstanding_reqs_i]);
				assign rdata_pmp_err_n[g_outstanding_reqs_i] = ((((valid_req & ~rdata_outstanding_q[g_outstanding_reqs_i]) & instr_pmp_err_i) & rdata_outstanding_q[(g_outstanding_reqs_i - 1)]) | rdata_pmp_err_q[g_outstanding_reqs_i]);
			end
		end
	endgenerate
	assign rdata_outstanding_s = (rvalid_or_pmp_err ? {1'b0, rdata_outstanding_n[(NUM_REQS - 1):1]} : rdata_outstanding_n);
	assign branch_discard_s = (rvalid_or_pmp_err ? {1'b0, branch_discard_n[(NUM_REQS - 1):1]} : branch_discard_n);
	assign rdata_pmp_err_s = (rvalid_or_pmp_err ? {1'b0, rdata_pmp_err_n[(NUM_REQS - 1):1]} : rdata_pmp_err_n);
	assign fifo_valid = (rvalid_or_pmp_err & ~branch_discard_q[0]);
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			valid_req_q <= 1'b0;
			discard_req_q <= 1'b0;
			rdata_outstanding_q <= 'b0;
			branch_discard_q <= 'b0;
			rdata_pmp_err_q <= 'b0;
		end
		else begin
			valid_req_q <= valid_req_d;
			discard_req_q <= discard_req_d;
			rdata_outstanding_q <= rdata_outstanding_s;
			branch_discard_q <= branch_discard_s;
			rdata_pmp_err_q <= rdata_pmp_err_s;
		end
	assign instr_req_o = valid_req;
	assign instr_addr_o = instr_addr_w_aligned;
endmodule
